


module sendblock();
	
	
	
endmodule
