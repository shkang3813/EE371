// Copyright (C) 2017  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel MegaCore Function License Agreement, or other 
// applicable license agreement, including, without limitation, 
// that your use is for the sole purpose of programming logic 
// devices manufactured by Intel and sold by Intel or its 
// authorized distributors.  Please refer to the applicable 
// agreement for further details.

// VENDOR "Altera"
// PROGRAM "Quartus Prime"
// VERSION "Version 17.0.2 Build 602 07/19/2017 SJ Standard Edition"

// DATE "12/05/2017 18:44:13"

// 
// Device: Altera 5CSEMA5F31C6 Package FBGA896
// 

// 
// This greybox netlist file is for third party Synthesis Tools
// for timing and resource estimation only.
// 


module first_nios2_system (
	altera_reserved_tms,
	altera_reserved_tck,
	altera_reserved_tdi,
	altera_reserved_tdo,
	camdata1_external_connection_export,
	camdata2_external_connection_export,
	camstate1_external_connection_export,
	camstate2_external_connection_export,
	clk_clk,
	download1_external_connection_export,
	download2_external_connection_export,
	hex1_external_connection_export,
	hex2_external_connection_export,
	leds_external_connection_export,
	reset_reset_n,
	rtd1_external_connection_export,
	rtd2_external_connection_export,
	start_external_connection_export,
	tenout1_external_connection_export,
	tenout2_external_connection_export)/* synthesis synthesis_greybox=1 */;
input 	altera_reserved_tms;
input 	altera_reserved_tck;
input 	altera_reserved_tdi;
output 	altera_reserved_tdo;
input 	[6:0] camdata1_external_connection_export;
input 	[6:0] camdata2_external_connection_export;
input 	[5:0] camstate1_external_connection_export;
input 	[5:0] camstate2_external_connection_export;
input 	clk_clk;
output 	download1_external_connection_export;
output 	download2_external_connection_export;
output 	[6:0] hex1_external_connection_export;
output 	[6:0] hex2_external_connection_export;
output 	[7:0] leds_external_connection_export;
input 	reset_reset_n;
input 	rtd1_external_connection_export;
input 	rtd2_external_connection_export;
output 	start_external_connection_export;
input 	[3:0] tenout1_external_connection_export;
input 	[3:0] tenout2_external_connection_export;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \onchip_mem|the_altsyncram|auto_generated|q_a[0] ;
wire \onchip_mem|the_altsyncram|auto_generated|q_a[1] ;
wire \onchip_mem|the_altsyncram|auto_generated|q_a[2] ;
wire \onchip_mem|the_altsyncram|auto_generated|q_a[3] ;
wire \onchip_mem|the_altsyncram|auto_generated|q_a[4] ;
wire \onchip_mem|the_altsyncram|auto_generated|q_a[5] ;
wire \onchip_mem|the_altsyncram|auto_generated|q_a[6] ;
wire \onchip_mem|the_altsyncram|auto_generated|q_a[7] ;
wire \mm_interconnect_0|jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[22]~q ;
wire \onchip_mem|the_altsyncram|auto_generated|q_a[22] ;
wire \onchip_mem|the_altsyncram|auto_generated|q_a[23] ;
wire \onchip_mem|the_altsyncram|auto_generated|q_a[24] ;
wire \onchip_mem|the_altsyncram|auto_generated|q_a[25] ;
wire \onchip_mem|the_altsyncram|auto_generated|q_a[31] ;
wire \onchip_mem|the_altsyncram|auto_generated|q_a[21] ;
wire \onchip_mem|the_altsyncram|auto_generated|q_a[11] ;
wire \onchip_mem|the_altsyncram|auto_generated|q_a[28] ;
wire \onchip_mem|the_altsyncram|auto_generated|q_a[10] ;
wire \onchip_mem|the_altsyncram|auto_generated|q_a[27] ;
wire \onchip_mem|the_altsyncram|auto_generated|q_a[8] ;
wire \onchip_mem|the_altsyncram|auto_generated|q_a[9] ;
wire \onchip_mem|the_altsyncram|auto_generated|q_a[26] ;
wire \mm_interconnect_0|jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[20]~q ;
wire \onchip_mem|the_altsyncram|auto_generated|q_a[20] ;
wire \mm_interconnect_0|jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[19]~q ;
wire \onchip_mem|the_altsyncram|auto_generated|q_a[19] ;
wire \onchip_mem|the_altsyncram|auto_generated|q_a[17] ;
wire \onchip_mem|the_altsyncram|auto_generated|q_a[30] ;
wire \onchip_mem|the_altsyncram|auto_generated|q_a[18] ;
wire \onchip_mem|the_altsyncram|auto_generated|q_a[16] ;
wire \onchip_mem|the_altsyncram|auto_generated|q_a[15] ;
wire \onchip_mem|the_altsyncram|auto_generated|q_a[12] ;
wire \onchip_mem|the_altsyncram|auto_generated|q_a[13] ;
wire \onchip_mem|the_altsyncram|auto_generated|q_a[14] ;
wire \onchip_mem|the_altsyncram|auto_generated|q_a[29] ;
wire \cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[0]~q ;
wire \camstate2|readdata[0]~q ;
wire \tenout1|readdata[0]~q ;
wire \tenout2|readdata[0]~q ;
wire \camstate1|readdata[0]~q ;
wire \rtd2|readdata[0]~q ;
wire \rtd1|readdata[0]~q ;
wire \jtag_uart|the_first_nios2_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[0] ;
wire \camdata1|readdata[0]~q ;
wire \camdata2|readdata[0]~q ;
wire \tenout2|readdata[1]~q ;
wire \cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[1]~q ;
wire \camdata1|readdata[1]~q ;
wire \camstate2|readdata[1]~q ;
wire \jtag_uart|the_first_nios2_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[1] ;
wire \camdata2|readdata[1]~q ;
wire \camstate1|readdata[1]~q ;
wire \tenout1|readdata[1]~q ;
wire \tenout2|readdata[2]~q ;
wire \cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[2]~q ;
wire \camdata1|readdata[2]~q ;
wire \camstate2|readdata[2]~q ;
wire \jtag_uart|the_first_nios2_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[2] ;
wire \camdata2|readdata[2]~q ;
wire \camstate1|readdata[2]~q ;
wire \tenout1|readdata[2]~q ;
wire \camdata2|readdata[3]~q ;
wire \tenout2|readdata[3]~q ;
wire \cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[3]~q ;
wire \camdata1|readdata[3]~q ;
wire \tenout1|readdata[3]~q ;
wire \jtag_uart|the_first_nios2_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[3] ;
wire \camstate1|readdata[3]~q ;
wire \camstate2|readdata[3]~q ;
wire \jtag_uart|the_first_nios2_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[4] ;
wire \cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[4]~q ;
wire \camdata1|readdata[4]~q ;
wire \camdata2|readdata[4]~q ;
wire \camstate1|readdata[4]~q ;
wire \camstate2|readdata[4]~q ;
wire \cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[5]~q ;
wire \camdata1|readdata[5]~q ;
wire \camdata2|readdata[5]~q ;
wire \jtag_uart|the_first_nios2_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[5] ;
wire \camstate1|readdata[5]~q ;
wire \camstate2|readdata[5]~q ;
wire \camdata1|readdata[6]~q ;
wire \jtag_uart|the_first_nios2_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[6] ;
wire \cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[6]~q ;
wire \camdata2|readdata[6]~q ;
wire \jtag_uart|the_first_nios2_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[7] ;
wire \cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[7]~q ;
wire \jtag_uart|Add1~1_sumout ;
wire \cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[22]~q ;
wire \cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[23]~q ;
wire \cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[24]~q ;
wire \cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[25]~q ;
wire \cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[31]~q ;
wire \cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[21]~q ;
wire \jtag_uart|Add1~5_sumout ;
wire \cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[11]~q ;
wire \cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[28]~q ;
wire \cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[10]~q ;
wire \cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[27]~q ;
wire \cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[8]~q ;
wire \cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[9]~q ;
wire \cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[26]~q ;
wire \jtag_uart|Add1~9_sumout ;
wire \cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[20]~q ;
wire \jtag_uart|Add1~13_sumout ;
wire \cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[19]~q ;
wire \cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[17]~q ;
wire \jtag_uart|Add1~17_sumout ;
wire \cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[30]~q ;
wire \cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[18]~q ;
wire \jtag_uart|Add1~21_sumout ;
wire \cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[16]~q ;
wire \jtag_uart|Add1~25_sumout ;
wire \cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[15]~q ;
wire \cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[12]~q ;
wire \cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[13]~q ;
wire \cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[14]~q ;
wire \cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[29]~q ;
wire \download1|data_out~q ;
wire \download2|data_out~q ;
wire \hex1|data_out[0]~q ;
wire \hex1|data_out[1]~q ;
wire \hex1|data_out[2]~q ;
wire \hex1|data_out[3]~q ;
wire \hex1|data_out[4]~q ;
wire \hex1|data_out[5]~q ;
wire \hex1|data_out[6]~q ;
wire \hex2|data_out[0]~q ;
wire \hex2|data_out[1]~q ;
wire \hex2|data_out[2]~q ;
wire \hex2|data_out[3]~q ;
wire \hex2|data_out[4]~q ;
wire \hex2|data_out[5]~q ;
wire \hex2|data_out[6]~q ;
wire \leds|data_out[0]~q ;
wire \leds|data_out[1]~q ;
wire \leds|data_out[2]~q ;
wire \leds|data_out[3]~q ;
wire \leds|data_out[4]~q ;
wire \leds|data_out[5]~q ;
wire \leds|data_out[6]~q ;
wire \leds|data_out[7]~q ;
wire \start|data_out~q ;
wire \cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[0]~q ;
wire \cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_tck|ir_out[0]~q ;
wire \cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_tck|ir_out[1]~q ;
wire \jtag_uart|first_nios2_system_jtag_uart_alt_jtag_atlantic|tdo~q ;
wire \cpu|cpu|A_st_data[0]~q ;
wire \mm_interconnect_0|download1_s1_agent_rsp_fifo|mem_used[1]~q ;
wire \cpu|cpu|A_mem_baddr[4]~q ;
wire \cpu|cpu|A_mem_baddr[5]~q ;
wire \cpu|cpu|A_mem_baddr[8]~q ;
wire \cpu|cpu|A_mem_baddr[16]~q ;
wire \cpu|cpu|A_mem_baddr[15]~q ;
wire \cpu|cpu|A_mem_baddr[14]~q ;
wire \cpu|cpu|A_mem_baddr[13]~q ;
wire \mm_interconnect_0|router|Equal1~0_combout ;
wire \cpu|cpu|A_mem_baddr[12]~q ;
wire \cpu|cpu|A_mem_baddr[11]~q ;
wire \cpu|cpu|A_mem_baddr[10]~q ;
wire \cpu|cpu|A_mem_baddr[9]~q ;
wire \mm_interconnect_0|router|Equal2~0_combout ;
wire \cpu|cpu|A_mem_baddr[7]~q ;
wire \cpu|cpu|A_mem_baddr[6]~q ;
wire \mm_interconnect_0|router|Equal15~1_combout ;
wire \download1|always0~0_combout ;
wire \cpu|cpu|clr_break_line~q ;
wire \mm_interconnect_0|download1_s1_translator|wait_latency_counter[1]~q ;
wire \mm_interconnect_0|download1_s1_translator|wait_latency_counter[0]~q ;
wire \cpu|cpu|d_write~q ;
wire \cpu|cpu|A_mem_baddr[3]~q ;
wire \cpu|cpu|A_mem_baddr[2]~q ;
wire \camdata1|Equal0~0_combout ;
wire \rst_controller|r_sync_rst~q ;
wire \mm_interconnect_0|download2_s1_agent_rsp_fifo|write~0_combout ;
wire \mm_interconnect_0|download2_s1_translator|wait_latency_counter[0]~q ;
wire \mm_interconnect_0|hex1_s1_translator|wait_latency_counter[1]~q ;
wire \mm_interconnect_0|hex1_s1_agent_rsp_fifo|mem_used[1]~q ;
wire \mm_interconnect_0|router|Equal6~1_combout ;
wire \mm_interconnect_0|hex1_s1_translator|wait_latency_counter[0]~q ;
wire \cpu|cpu|A_st_data[1]~q ;
wire \cpu|cpu|A_st_data[2]~q ;
wire \cpu|cpu|A_st_data[3]~q ;
wire \cpu|cpu|A_st_data[4]~q ;
wire \cpu|cpu|A_st_data[5]~q ;
wire \cpu|cpu|A_st_data[6]~q ;
wire \mm_interconnect_0|hex2_s1_translator|wait_latency_counter[1]~q ;
wire \mm_interconnect_0|hex2_s1_agent_rsp_fifo|mem_used[1]~q ;
wire \mm_interconnect_0|router|always1~0_combout ;
wire \mm_interconnect_0|hex2_s1_translator|wait_latency_counter[0]~q ;
wire \mm_interconnect_0|leds_s1_translator|wait_latency_counter[1]~q ;
wire \mm_interconnect_0|leds_s1_agent_rsp_fifo|mem_used[1]~q ;
wire \mm_interconnect_0|router|Equal16~0_combout ;
wire \mm_interconnect_0|leds_s1_translator|wait_latency_counter[0]~q ;
wire \cpu|cpu|A_st_data[7]~q ;
wire \mm_interconnect_0|start_s1_translator|wait_latency_counter[1]~q ;
wire \mm_interconnect_0|start_s1_agent|m0_write~0_combout ;
wire \mm_interconnect_0|start_s1_translator|wait_latency_counter[0]~q ;
wire \cpu|cpu|d_read~q ;
wire \mm_interconnect_0|download1_s1_translator|read_latency_shift_reg~0_combout ;
wire \mm_interconnect_0|cpu_data_master_agent|cp_valid~0_combout ;
wire \cpu|cpu|W_debug_mode~q ;
wire \mm_interconnect_0|camstate1_s1_translator|read_latency_shift_reg[0]~q ;
wire \mm_interconnect_0|rsp_mux|WideOr1~0_combout ;
wire \mm_interconnect_0|rsp_mux|WideOr1~1_combout ;
wire \mm_interconnect_0|rsp_demux_002|src0_valid~0_combout ;
wire \mm_interconnect_0|rsp_demux_003|src0_valid~0_combout ;
wire \mm_interconnect_0|jtag_uart_avalon_jtag_slave_translator|read_latency_shift_reg[0]~q ;
wire \mm_interconnect_0|rsp_mux|WideOr1~3_combout ;
wire \mm_interconnect_0|rsp_mux|WideOr1~combout ;
wire \mm_interconnect_0|router|Equal2~2_combout ;
wire \mm_interconnect_0|sys_clk_timer_s1_translator|wait_latency_counter[0]~q ;
wire \mm_interconnect_0|sys_clk_timer_s1_agent_rsp_fifo|mem_used[1]~q ;
wire \mm_interconnect_0|sys_clk_timer_s1_translator|wait_latency_counter[1]~q ;
wire \mm_interconnect_0|onchip_mem_s1_agent_rsp_fifo|mem_used[1]~q ;
wire \mm_interconnect_0|cmd_mux_003|saved_grant[0]~q ;
wire \mm_interconnect_0|router|always1~2_combout ;
wire \jtag_uart|av_waitrequest~q ;
wire \mm_interconnect_0|jtag_uart_avalon_jtag_slave_agent_rsp_fifo|mem_used[1]~q ;
wire \jtag_uart|av_waitrequest~0_combout ;
wire \mm_interconnect_0|cmd_mux_002|saved_grant[0]~q ;
wire \cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|the_first_nios2_system_cpu_cpu_nios2_ocimem|waitrequest~q ;
wire \mm_interconnect_0|cpu_debug_mem_slave_agent_rsp_fifo|mem_used[1]~q ;
wire \mm_interconnect_0|cpu_data_master_translator|av_waitrequest~0_combout ;
wire \cpu|cpu|i_read~q ;
wire \cpu|cpu|ic_fill_tag[5]~q ;
wire \cpu|cpu|ic_fill_tag[4]~q ;
wire \cpu|cpu|ic_fill_tag[3]~q ;
wire \cpu|cpu|ic_fill_tag[2]~q ;
wire \cpu|cpu|ic_fill_tag[1]~q ;
wire \cpu|cpu|ic_fill_tag[0]~q ;
wire \mm_interconnect_0|cmd_mux_002|WideOr1~combout ;
wire \mm_interconnect_0|cpu_debug_mem_slave_agent_rsp_fifo|mem~0_combout ;
wire \mm_interconnect_0|cmd_mux_003|WideOr1~combout ;
wire \sys_clk_timer|timeout_occurred~q ;
wire \sys_clk_timer|control_register[0]~q ;
wire \jtag_uart|ien_AE~q ;
wire \jtag_uart|av_readdata[9]~combout ;
wire \jtag_uart|ien_AF~q ;
wire \jtag_uart|av_readdata[8]~0_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~0_combout ;
wire \cpu|cpu|ic_fill_ap_offset[0]~q ;
wire \mm_interconnect_0|cmd_mux_002|src_data[38]~combout ;
wire \cpu|cpu|ic_fill_line[0]~q ;
wire \mm_interconnect_0|cmd_mux_002|src_data[41]~combout ;
wire \cpu|cpu|ic_fill_ap_offset[2]~q ;
wire \mm_interconnect_0|cmd_mux_002|src_data[40]~combout ;
wire \cpu|cpu|ic_fill_ap_offset[1]~q ;
wire \mm_interconnect_0|cmd_mux_002|src_data[39]~combout ;
wire \cpu|cpu|ic_fill_line[5]~q ;
wire \mm_interconnect_0|cmd_mux_002|src_data[46]~combout ;
wire \cpu|cpu|ic_fill_line[4]~q ;
wire \mm_interconnect_0|cmd_mux_002|src_data[45]~combout ;
wire \cpu|cpu|ic_fill_line[3]~q ;
wire \mm_interconnect_0|cmd_mux_002|src_data[44]~combout ;
wire \cpu|cpu|ic_fill_line[2]~q ;
wire \mm_interconnect_0|cmd_mux_002|src_data[43]~combout ;
wire \cpu|cpu|ic_fill_line[1]~q ;
wire \mm_interconnect_0|cmd_mux_002|src_data[42]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~1_combout ;
wire \mm_interconnect_0|cpu_instruction_master_limiter|save_dest_id~0_combout ;
wire \mm_interconnect_0|cmd_demux_001|WideOr0~0_combout ;
wire \mm_interconnect_0|cpu_instruction_master_limiter|nonposted_cmd_accepted~combout ;
wire \mm_interconnect_0|cpu_instruction_master_limiter|suppress_change_dest_id~0_combout ;
wire \rst_controller|r_early_rst~q ;
wire \jtag_uart|the_first_nios2_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|b_full~q ;
wire \mm_interconnect_0|rsp_mux|src_data[0]~combout ;
wire \jtag_uart|the_first_nios2_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|b_full~q ;
wire \jtag_uart|the_first_nios2_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|b_non_empty~q ;
wire \jtag_uart|read_0~q ;
wire \jtag_uart|the_first_nios2_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[0]~q ;
wire \mm_interconnect_0|rsp_mux|src_payload~0_combout ;
wire \mm_interconnect_0|rsp_mux|src_data[1]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[2]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[3]~combout ;
wire \mm_interconnect_0|rsp_mux|src_payload~3_combout ;
wire \mm_interconnect_0|rsp_mux|src_payload~7_combout ;
wire \mm_interconnect_0|rsp_mux|src_payload~12_combout ;
wire \mm_interconnect_0|rsp_mux|src_payload~15_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~2_combout ;
wire \cpu|cpu|A_mem_byte_en[0]~q ;
wire \mm_interconnect_0|cmd_mux_002|src_data[32]~combout ;
wire \jtag_uart|the_first_nios2_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[1]~q ;
wire \jtag_uart|the_first_nios2_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[4]~q ;
wire \jtag_uart|the_first_nios2_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[3]~q ;
wire \jtag_uart|the_first_nios2_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[2]~q ;
wire \jtag_uart|the_first_nios2_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[5]~q ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[22]~q ;
wire \mm_interconnect_0|rsp_mux|src_payload~16_combout ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[23]~q ;
wire \mm_interconnect_0|rsp_mux|src_payload~17_combout ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[24]~q ;
wire \mm_interconnect_0|rsp_mux|src_payload~18_combout ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[25]~q ;
wire \mm_interconnect_0|rsp_mux|src_payload~19_combout ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[31]~q ;
wire \mm_interconnect_0|rsp_mux|src_payload~20_combout ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[21]~q ;
wire \mm_interconnect_0|rsp_mux|src_payload~21_combout ;
wire \mm_interconnect_0|rsp_mux|src_payload~22_combout ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[11]~q ;
wire \mm_interconnect_0|rsp_mux|src_payload~23_combout ;
wire \mm_interconnect_0|rsp_mux|src_payload~24_combout ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[28]~q ;
wire \mm_interconnect_0|rsp_mux|src_payload~25_combout ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[10]~q ;
wire \mm_interconnect_0|rsp_mux|src_payload~26_combout ;
wire \mm_interconnect_0|rsp_mux|src_payload~27_combout ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[27]~q ;
wire \mm_interconnect_0|rsp_mux|src_payload~28_combout ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[8]~q ;
wire \mm_interconnect_0|rsp_mux|src_payload~29_combout ;
wire \mm_interconnect_0|rsp_mux|src_payload~30_combout ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[9]~q ;
wire \mm_interconnect_0|rsp_mux|src_payload~31_combout ;
wire \mm_interconnect_0|rsp_mux|src_payload~32_combout ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[26]~q ;
wire \mm_interconnect_0|rsp_mux|src_payload~33_combout ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[20]~q ;
wire \mm_interconnect_0|rsp_mux|src_payload~34_combout ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[19]~q ;
wire \mm_interconnect_0|rsp_mux|src_payload~35_combout ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[17]~q ;
wire \mm_interconnect_0|rsp_mux|src_payload~36_combout ;
wire \mm_interconnect_0|rsp_mux|src_payload~37_combout ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[30]~q ;
wire \mm_interconnect_0|rsp_mux|src_payload~38_combout ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[18]~q ;
wire \mm_interconnect_0|rsp_mux|src_payload~39_combout ;
wire \mm_interconnect_0|rsp_mux|src_payload~40_combout ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[16]~q ;
wire \mm_interconnect_0|rsp_mux|src_payload~41_combout ;
wire \mm_interconnect_0|rsp_mux|src_payload~42_combout ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[15]~q ;
wire \mm_interconnect_0|rsp_mux|src_payload~43_combout ;
wire \mm_interconnect_0|rsp_mux|src_payload~44_combout ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[12]~q ;
wire \mm_interconnect_0|rsp_mux|src_payload~45_combout ;
wire \mm_interconnect_0|rsp_mux|src_payload~46_combout ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[13]~q ;
wire \mm_interconnect_0|rsp_mux|src_payload~47_combout ;
wire \mm_interconnect_0|rsp_mux|src_payload~48_combout ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[14]~q ;
wire \mm_interconnect_0|rsp_mux|src_payload~49_combout ;
wire \mm_interconnect_0|rsp_mux|src_payload~50_combout ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[29]~q ;
wire \mm_interconnect_0|rsp_mux|src_payload~51_combout ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~0_combout ;
wire \mm_interconnect_0|cmd_mux_003|src_data[38]~combout ;
wire \mm_interconnect_0|cmd_mux_003|src_data[39]~combout ;
wire \mm_interconnect_0|cmd_mux_003|src_data[40]~combout ;
wire \mm_interconnect_0|cmd_mux_003|src_data[41]~combout ;
wire \mm_interconnect_0|cmd_mux_003|src_data[42]~combout ;
wire \mm_interconnect_0|cmd_mux_003|src_data[43]~combout ;
wire \mm_interconnect_0|cmd_mux_003|src_data[44]~combout ;
wire \mm_interconnect_0|cmd_mux_003|src_data[45]~combout ;
wire \mm_interconnect_0|cmd_mux_003|src_data[46]~combout ;
wire \mm_interconnect_0|cmd_mux_003|src_data[47]~combout ;
wire \mm_interconnect_0|cmd_mux_003|src_data[48]~combout ;
wire \mm_interconnect_0|cmd_mux_003|src_data[49]~combout ;
wire \mm_interconnect_0|cmd_mux_003|src_data[50]~combout ;
wire \mm_interconnect_0|cmd_mux_003|src_data[32]~combout ;
wire \sys_clk_timer|readdata[0]~q ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~3_combout ;
wire \cpu|cpu|A_st_data[16]~q ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~4_combout ;
wire \mm_interconnect_0|rsp_mux_001|WideOr1~combout ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~1_combout ;
wire \sys_clk_timer|readdata[1]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~2_combout ;
wire \sys_clk_timer|readdata[2]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~3_combout ;
wire \sys_clk_timer|readdata[3]~q ;
wire \sys_clk_timer|readdata[4]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~4_combout ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~5_combout ;
wire \sys_clk_timer|readdata[5]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~6_combout ;
wire \sys_clk_timer|readdata[6]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~7_combout ;
wire \sys_clk_timer|readdata[7]~q ;
wire \cpu|cpu|A_st_data[22]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~8_combout ;
wire \cpu|cpu|A_mem_byte_en[2]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_data[34]~combout ;
wire \cpu|cpu|A_st_data[23]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~9_combout ;
wire \cpu|cpu|A_st_data[24]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~10_combout ;
wire \cpu|cpu|A_mem_byte_en[3]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_data[35]~combout ;
wire \cpu|cpu|A_st_data[25]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~11_combout ;
wire \cpu|cpu|A_st_data[31]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~12_combout ;
wire \cpu|cpu|A_st_data[21]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~13_combout ;
wire \cpu|cpu|A_st_data[11]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~14_combout ;
wire \cpu|cpu|A_mem_byte_en[1]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_data[33]~combout ;
wire \sys_clk_timer|readdata[11]~q ;
wire \cpu|cpu|A_st_data[28]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~15_combout ;
wire \cpu|cpu|A_st_data[10]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~16_combout ;
wire \jtag_uart|ac~q ;
wire \sys_clk_timer|readdata[10]~q ;
wire \cpu|cpu|A_st_data[27]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~17_combout ;
wire \cpu|cpu|A_st_data[8]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~18_combout ;
wire \sys_clk_timer|readdata[8]~q ;
wire \cpu|cpu|A_st_data[9]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~19_combout ;
wire \sys_clk_timer|readdata[9]~q ;
wire \cpu|cpu|A_st_data[26]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~20_combout ;
wire \cpu|cpu|A_st_data[20]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~21_combout ;
wire \cpu|cpu|A_st_data[19]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~22_combout ;
wire \cpu|cpu|A_st_data[17]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~23_combout ;
wire \cpu|cpu|A_st_data[30]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~24_combout ;
wire \cpu|cpu|A_st_data[18]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~25_combout ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~26_combout ;
wire \cpu|cpu|A_st_data[15]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~27_combout ;
wire \jtag_uart|rvalid~q ;
wire \sys_clk_timer|readdata[15]~q ;
wire \cpu|cpu|A_st_data[12]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~28_combout ;
wire \sys_clk_timer|readdata[12]~q ;
wire \cpu|cpu|A_st_data[13]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~29_combout ;
wire \sys_clk_timer|readdata[13]~q ;
wire \cpu|cpu|A_st_data[14]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~30_combout ;
wire \jtag_uart|woverflow~q ;
wire \sys_clk_timer|readdata[14]~q ;
wire \cpu|cpu|A_st_data[29]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~31_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[26]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[25]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[24]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[23]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[22]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[1]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[0]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[2]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[3]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[4]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[5]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[28]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[31]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[27]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[29]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[30]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[11]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[12]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[13]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[14]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[15]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[16]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~5_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[9]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[21]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[6]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[8]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[17]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[18]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[10]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[7]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[20]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[19]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~6_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[34]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~7_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~8_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~9_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~10_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~11_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~12_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~13_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~14_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~15_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[35]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~16_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~17_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~18_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~19_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~20_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~21_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~22_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[33]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~23_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~24_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~25_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~26_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~27_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~28_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~29_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~30_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~31_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~32_combout ;
wire \rst_controller|alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain[1]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_1[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~14_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~7_combout ;
wire \auto_hub|~GND~combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell_combout ;
wire \clk_clk~input_o ;
wire \camstate2_external_connection_export[0]~input_o ;
wire \tenout1_external_connection_export[0]~input_o ;
wire \tenout2_external_connection_export[0]~input_o ;
wire \camstate1_external_connection_export[0]~input_o ;
wire \rtd2_external_connection_export~input_o ;
wire \rtd1_external_connection_export~input_o ;
wire \camdata1_external_connection_export[0]~input_o ;
wire \camdata2_external_connection_export[0]~input_o ;
wire \reset_reset_n~input_o ;
wire \tenout2_external_connection_export[1]~input_o ;
wire \camdata1_external_connection_export[1]~input_o ;
wire \camstate2_external_connection_export[1]~input_o ;
wire \camdata2_external_connection_export[1]~input_o ;
wire \camstate1_external_connection_export[1]~input_o ;
wire \tenout1_external_connection_export[1]~input_o ;
wire \tenout2_external_connection_export[2]~input_o ;
wire \camdata1_external_connection_export[2]~input_o ;
wire \camstate2_external_connection_export[2]~input_o ;
wire \camdata2_external_connection_export[2]~input_o ;
wire \camstate1_external_connection_export[2]~input_o ;
wire \tenout1_external_connection_export[2]~input_o ;
wire \camdata2_external_connection_export[3]~input_o ;
wire \tenout2_external_connection_export[3]~input_o ;
wire \camdata1_external_connection_export[3]~input_o ;
wire \tenout1_external_connection_export[3]~input_o ;
wire \camstate1_external_connection_export[3]~input_o ;
wire \camstate2_external_connection_export[3]~input_o ;
wire \camdata1_external_connection_export[4]~input_o ;
wire \camdata2_external_connection_export[4]~input_o ;
wire \camstate1_external_connection_export[4]~input_o ;
wire \camstate2_external_connection_export[4]~input_o ;
wire \camdata1_external_connection_export[5]~input_o ;
wire \camdata2_external_connection_export[5]~input_o ;
wire \camstate1_external_connection_export[5]~input_o ;
wire \camstate2_external_connection_export[5]~input_o ;
wire \camdata1_external_connection_export[6]~input_o ;
wire \camdata2_external_connection_export[6]~input_o ;
wire \altera_reserved_tms~input_o ;
wire \altera_reserved_tck~input_o ;
wire \altera_reserved_tdi~input_o ;
wire \altera_internal_jtag~TCKUTAP ;
wire \altera_internal_jtag~TMSUTAP ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ;
wire \altera_internal_jtag~TDIUTAP ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ;
wire \~GND~combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~8_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~10_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~q ;
wire \altera_internal_jtag~TDO ;


first_nios2_system_first_nios2_system_cpu cpu(
	.av_readdata_pre_22(\mm_interconnect_0|jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[22]~q ),
	.q_a_22(\onchip_mem|the_altsyncram|auto_generated|q_a[22] ),
	.q_a_23(\onchip_mem|the_altsyncram|auto_generated|q_a[23] ),
	.q_a_24(\onchip_mem|the_altsyncram|auto_generated|q_a[24] ),
	.q_a_25(\onchip_mem|the_altsyncram|auto_generated|q_a[25] ),
	.q_a_31(\onchip_mem|the_altsyncram|auto_generated|q_a[31] ),
	.q_a_21(\onchip_mem|the_altsyncram|auto_generated|q_a[21] ),
	.q_a_11(\onchip_mem|the_altsyncram|auto_generated|q_a[11] ),
	.q_a_28(\onchip_mem|the_altsyncram|auto_generated|q_a[28] ),
	.q_a_10(\onchip_mem|the_altsyncram|auto_generated|q_a[10] ),
	.q_a_27(\onchip_mem|the_altsyncram|auto_generated|q_a[27] ),
	.q_a_8(\onchip_mem|the_altsyncram|auto_generated|q_a[8] ),
	.q_a_9(\onchip_mem|the_altsyncram|auto_generated|q_a[9] ),
	.q_a_26(\onchip_mem|the_altsyncram|auto_generated|q_a[26] ),
	.av_readdata_pre_20(\mm_interconnect_0|jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[20]~q ),
	.q_a_20(\onchip_mem|the_altsyncram|auto_generated|q_a[20] ),
	.av_readdata_pre_19(\mm_interconnect_0|jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[19]~q ),
	.q_a_19(\onchip_mem|the_altsyncram|auto_generated|q_a[19] ),
	.q_a_17(\onchip_mem|the_altsyncram|auto_generated|q_a[17] ),
	.q_a_30(\onchip_mem|the_altsyncram|auto_generated|q_a[30] ),
	.q_a_18(\onchip_mem|the_altsyncram|auto_generated|q_a[18] ),
	.q_a_16(\onchip_mem|the_altsyncram|auto_generated|q_a[16] ),
	.q_a_15(\onchip_mem|the_altsyncram|auto_generated|q_a[15] ),
	.q_a_12(\onchip_mem|the_altsyncram|auto_generated|q_a[12] ),
	.q_a_13(\onchip_mem|the_altsyncram|auto_generated|q_a[13] ),
	.q_a_14(\onchip_mem|the_altsyncram|auto_generated|q_a[14] ),
	.q_a_29(\onchip_mem|the_altsyncram|auto_generated|q_a[29] ),
	.readdata_0(\cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[0]~q ),
	.readdata_1(\cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[1]~q ),
	.readdata_2(\cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[2]~q ),
	.readdata_3(\cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[3]~q ),
	.readdata_4(\cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[4]~q ),
	.readdata_5(\cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[5]~q ),
	.readdata_6(\cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[6]~q ),
	.readdata_7(\cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[7]~q ),
	.readdata_22(\cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[22]~q ),
	.readdata_23(\cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[23]~q ),
	.readdata_24(\cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[24]~q ),
	.readdata_25(\cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[25]~q ),
	.readdata_31(\cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[31]~q ),
	.readdata_21(\cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[21]~q ),
	.readdata_11(\cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[11]~q ),
	.readdata_28(\cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[28]~q ),
	.readdata_10(\cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[10]~q ),
	.readdata_27(\cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[27]~q ),
	.readdata_8(\cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[8]~q ),
	.readdata_9(\cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[9]~q ),
	.readdata_26(\cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[26]~q ),
	.readdata_20(\cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[20]~q ),
	.readdata_19(\cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[19]~q ),
	.readdata_17(\cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[17]~q ),
	.readdata_30(\cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[30]~q ),
	.readdata_18(\cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[18]~q ),
	.readdata_16(\cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[16]~q ),
	.readdata_15(\cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[15]~q ),
	.readdata_12(\cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[12]~q ),
	.readdata_13(\cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[13]~q ),
	.readdata_14(\cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[14]~q ),
	.readdata_29(\cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[29]~q ),
	.sr_0(\cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[0]~q ),
	.ir_out_0(\cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_tck|ir_out[0]~q ),
	.ir_out_1(\cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_tck|ir_out[1]~q ),
	.A_st_data_0(\cpu|cpu|A_st_data[0]~q ),
	.A_mem_baddr_4(\cpu|cpu|A_mem_baddr[4]~q ),
	.A_mem_baddr_5(\cpu|cpu|A_mem_baddr[5]~q ),
	.A_mem_baddr_8(\cpu|cpu|A_mem_baddr[8]~q ),
	.A_mem_baddr_16(\cpu|cpu|A_mem_baddr[16]~q ),
	.A_mem_baddr_15(\cpu|cpu|A_mem_baddr[15]~q ),
	.A_mem_baddr_14(\cpu|cpu|A_mem_baddr[14]~q ),
	.A_mem_baddr_13(\cpu|cpu|A_mem_baddr[13]~q ),
	.A_mem_baddr_12(\cpu|cpu|A_mem_baddr[12]~q ),
	.A_mem_baddr_11(\cpu|cpu|A_mem_baddr[11]~q ),
	.A_mem_baddr_10(\cpu|cpu|A_mem_baddr[10]~q ),
	.A_mem_baddr_9(\cpu|cpu|A_mem_baddr[9]~q ),
	.A_mem_baddr_7(\cpu|cpu|A_mem_baddr[7]~q ),
	.A_mem_baddr_6(\cpu|cpu|A_mem_baddr[6]~q ),
	.clr_break_line(\cpu|cpu|clr_break_line~q ),
	.d_write(\cpu|cpu|d_write~q ),
	.A_mem_baddr_3(\cpu|cpu|A_mem_baddr[3]~q ),
	.A_mem_baddr_2(\cpu|cpu|A_mem_baddr[2]~q ),
	.r_sync_rst(\rst_controller|r_sync_rst~q ),
	.A_st_data_1(\cpu|cpu|A_st_data[1]~q ),
	.A_st_data_2(\cpu|cpu|A_st_data[2]~q ),
	.A_st_data_3(\cpu|cpu|A_st_data[3]~q ),
	.A_st_data_4(\cpu|cpu|A_st_data[4]~q ),
	.A_st_data_5(\cpu|cpu|A_st_data[5]~q ),
	.A_st_data_6(\cpu|cpu|A_st_data[6]~q ),
	.A_st_data_7(\cpu|cpu|A_st_data[7]~q ),
	.d_read(\cpu|cpu|d_read~q ),
	.W_debug_mode(\cpu|cpu|W_debug_mode~q ),
	.read_latency_shift_reg_0(\mm_interconnect_0|camstate1_s1_translator|read_latency_shift_reg[0]~q ),
	.WideOr1(\mm_interconnect_0|rsp_mux|WideOr1~0_combout ),
	.WideOr11(\mm_interconnect_0|rsp_mux|WideOr1~1_combout ),
	.src0_valid(\mm_interconnect_0|rsp_demux_002|src0_valid~0_combout ),
	.src0_valid1(\mm_interconnect_0|rsp_demux_003|src0_valid~0_combout ),
	.read_latency_shift_reg_01(\mm_interconnect_0|jtag_uart_avalon_jtag_slave_translator|read_latency_shift_reg[0]~q ),
	.WideOr12(\mm_interconnect_0|rsp_mux|WideOr1~3_combout ),
	.WideOr13(\mm_interconnect_0|rsp_mux|WideOr1~combout ),
	.saved_grant_0(\mm_interconnect_0|cmd_mux_002|saved_grant[0]~q ),
	.debug_mem_slave_waitrequest(\cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|the_first_nios2_system_cpu_cpu_nios2_ocimem|waitrequest~q ),
	.mem_used_1(\mm_interconnect_0|cpu_debug_mem_slave_agent_rsp_fifo|mem_used[1]~q ),
	.av_waitrequest(\mm_interconnect_0|cpu_data_master_translator|av_waitrequest~0_combout ),
	.i_read(\cpu|cpu|i_read~q ),
	.ic_fill_tag_5(\cpu|cpu|ic_fill_tag[5]~q ),
	.ic_fill_tag_4(\cpu|cpu|ic_fill_tag[4]~q ),
	.ic_fill_tag_3(\cpu|cpu|ic_fill_tag[3]~q ),
	.ic_fill_tag_2(\cpu|cpu|ic_fill_tag[2]~q ),
	.ic_fill_tag_1(\cpu|cpu|ic_fill_tag[1]~q ),
	.ic_fill_tag_0(\cpu|cpu|ic_fill_tag[0]~q ),
	.WideOr14(\mm_interconnect_0|cmd_mux_002|WideOr1~combout ),
	.mem(\mm_interconnect_0|cpu_debug_mem_slave_agent_rsp_fifo|mem~0_combout ),
	.timeout_occurred(\sys_clk_timer|timeout_occurred~q ),
	.control_register_0(\sys_clk_timer|control_register[0]~q ),
	.av_readdata_9(\jtag_uart|av_readdata[9]~combout ),
	.av_readdata_8(\jtag_uart|av_readdata[8]~0_combout ),
	.src_payload(\mm_interconnect_0|cmd_mux_002|src_payload~0_combout ),
	.ic_fill_ap_offset_0(\cpu|cpu|ic_fill_ap_offset[0]~q ),
	.src_data_38(\mm_interconnect_0|cmd_mux_002|src_data[38]~combout ),
	.ic_fill_line_0(\cpu|cpu|ic_fill_line[0]~q ),
	.src_data_41(\mm_interconnect_0|cmd_mux_002|src_data[41]~combout ),
	.ic_fill_ap_offset_2(\cpu|cpu|ic_fill_ap_offset[2]~q ),
	.src_data_40(\mm_interconnect_0|cmd_mux_002|src_data[40]~combout ),
	.ic_fill_ap_offset_1(\cpu|cpu|ic_fill_ap_offset[1]~q ),
	.src_data_39(\mm_interconnect_0|cmd_mux_002|src_data[39]~combout ),
	.ic_fill_line_5(\cpu|cpu|ic_fill_line[5]~q ),
	.src_data_46(\mm_interconnect_0|cmd_mux_002|src_data[46]~combout ),
	.ic_fill_line_4(\cpu|cpu|ic_fill_line[4]~q ),
	.src_data_45(\mm_interconnect_0|cmd_mux_002|src_data[45]~combout ),
	.ic_fill_line_3(\cpu|cpu|ic_fill_line[3]~q ),
	.src_data_44(\mm_interconnect_0|cmd_mux_002|src_data[44]~combout ),
	.ic_fill_line_2(\cpu|cpu|ic_fill_line[2]~q ),
	.src_data_43(\mm_interconnect_0|cmd_mux_002|src_data[43]~combout ),
	.ic_fill_line_1(\cpu|cpu|ic_fill_line[1]~q ),
	.src_data_42(\mm_interconnect_0|cmd_mux_002|src_data[42]~combout ),
	.src_payload1(\mm_interconnect_0|cmd_mux_002|src_payload~1_combout ),
	.save_dest_id(\mm_interconnect_0|cpu_instruction_master_limiter|save_dest_id~0_combout ),
	.WideOr0(\mm_interconnect_0|cmd_demux_001|WideOr0~0_combout ),
	.nonposted_cmd_accepted(\mm_interconnect_0|cpu_instruction_master_limiter|nonposted_cmd_accepted~combout ),
	.suppress_change_dest_id(\mm_interconnect_0|cpu_instruction_master_limiter|suppress_change_dest_id~0_combout ),
	.r_early_rst(\rst_controller|r_early_rst~q ),
	.src_data_0(\mm_interconnect_0|rsp_mux|src_data[0]~combout ),
	.src_payload2(\mm_interconnect_0|rsp_mux|src_payload~0_combout ),
	.src_data_1(\mm_interconnect_0|rsp_mux|src_data[1]~combout ),
	.src_data_2(\mm_interconnect_0|rsp_mux|src_data[2]~combout ),
	.src_data_3(\mm_interconnect_0|rsp_mux|src_data[3]~combout ),
	.src_payload3(\mm_interconnect_0|rsp_mux|src_payload~3_combout ),
	.src_payload4(\mm_interconnect_0|rsp_mux|src_payload~7_combout ),
	.src_payload5(\mm_interconnect_0|rsp_mux|src_payload~12_combout ),
	.src_payload6(\mm_interconnect_0|rsp_mux|src_payload~15_combout ),
	.src_payload7(\mm_interconnect_0|cmd_mux_002|src_payload~2_combout ),
	.A_mem_byte_en_0(\cpu|cpu|A_mem_byte_en[0]~q ),
	.src_data_32(\mm_interconnect_0|cmd_mux_002|src_data[32]~combout ),
	.av_readdata_pre_221(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[22]~q ),
	.src_payload8(\mm_interconnect_0|rsp_mux|src_payload~16_combout ),
	.av_readdata_pre_23(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[23]~q ),
	.src_payload9(\mm_interconnect_0|rsp_mux|src_payload~17_combout ),
	.av_readdata_pre_24(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[24]~q ),
	.src_payload10(\mm_interconnect_0|rsp_mux|src_payload~18_combout ),
	.av_readdata_pre_25(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[25]~q ),
	.src_payload11(\mm_interconnect_0|rsp_mux|src_payload~19_combout ),
	.av_readdata_pre_31(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[31]~q ),
	.src_payload12(\mm_interconnect_0|rsp_mux|src_payload~20_combout ),
	.av_readdata_pre_21(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[21]~q ),
	.src_payload13(\mm_interconnect_0|rsp_mux|src_payload~21_combout ),
	.src_payload14(\mm_interconnect_0|rsp_mux|src_payload~22_combout ),
	.av_readdata_pre_11(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[11]~q ),
	.src_payload15(\mm_interconnect_0|rsp_mux|src_payload~23_combout ),
	.src_payload16(\mm_interconnect_0|rsp_mux|src_payload~24_combout ),
	.av_readdata_pre_28(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[28]~q ),
	.src_payload17(\mm_interconnect_0|rsp_mux|src_payload~25_combout ),
	.av_readdata_pre_10(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[10]~q ),
	.src_payload18(\mm_interconnect_0|rsp_mux|src_payload~26_combout ),
	.src_payload19(\mm_interconnect_0|rsp_mux|src_payload~27_combout ),
	.av_readdata_pre_27(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[27]~q ),
	.src_payload20(\mm_interconnect_0|rsp_mux|src_payload~28_combout ),
	.av_readdata_pre_8(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[8]~q ),
	.src_payload21(\mm_interconnect_0|rsp_mux|src_payload~29_combout ),
	.src_payload22(\mm_interconnect_0|rsp_mux|src_payload~30_combout ),
	.av_readdata_pre_9(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[9]~q ),
	.src_payload23(\mm_interconnect_0|rsp_mux|src_payload~31_combout ),
	.src_payload24(\mm_interconnect_0|rsp_mux|src_payload~32_combout ),
	.av_readdata_pre_26(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[26]~q ),
	.src_payload25(\mm_interconnect_0|rsp_mux|src_payload~33_combout ),
	.av_readdata_pre_201(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[20]~q ),
	.src_payload26(\mm_interconnect_0|rsp_mux|src_payload~34_combout ),
	.av_readdata_pre_191(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[19]~q ),
	.src_payload27(\mm_interconnect_0|rsp_mux|src_payload~35_combout ),
	.av_readdata_pre_17(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[17]~q ),
	.src_payload28(\mm_interconnect_0|rsp_mux|src_payload~36_combout ),
	.src_payload29(\mm_interconnect_0|rsp_mux|src_payload~37_combout ),
	.av_readdata_pre_30(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[30]~q ),
	.src_payload30(\mm_interconnect_0|rsp_mux|src_payload~38_combout ),
	.av_readdata_pre_18(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[18]~q ),
	.src_payload31(\mm_interconnect_0|rsp_mux|src_payload~39_combout ),
	.src_payload32(\mm_interconnect_0|rsp_mux|src_payload~40_combout ),
	.av_readdata_pre_16(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[16]~q ),
	.src_payload33(\mm_interconnect_0|rsp_mux|src_payload~41_combout ),
	.src_payload34(\mm_interconnect_0|rsp_mux|src_payload~42_combout ),
	.av_readdata_pre_15(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[15]~q ),
	.src_payload35(\mm_interconnect_0|rsp_mux|src_payload~43_combout ),
	.src_payload36(\mm_interconnect_0|rsp_mux|src_payload~44_combout ),
	.av_readdata_pre_12(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[12]~q ),
	.src_payload37(\mm_interconnect_0|rsp_mux|src_payload~45_combout ),
	.src_payload38(\mm_interconnect_0|rsp_mux|src_payload~46_combout ),
	.av_readdata_pre_13(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[13]~q ),
	.src_payload39(\mm_interconnect_0|rsp_mux|src_payload~47_combout ),
	.src_payload40(\mm_interconnect_0|rsp_mux|src_payload~48_combout ),
	.av_readdata_pre_14(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[14]~q ),
	.src_payload41(\mm_interconnect_0|rsp_mux|src_payload~49_combout ),
	.src_payload42(\mm_interconnect_0|rsp_mux|src_payload~50_combout ),
	.av_readdata_pre_29(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[29]~q ),
	.src_payload43(\mm_interconnect_0|rsp_mux|src_payload~51_combout ),
	.src_payload44(\mm_interconnect_0|cmd_mux_002|src_payload~3_combout ),
	.A_st_data_16(\cpu|cpu|A_st_data[16]~q ),
	.src_payload45(\mm_interconnect_0|cmd_mux_002|src_payload~4_combout ),
	.WideOr15(\mm_interconnect_0|rsp_mux_001|WideOr1~combout ),
	.A_st_data_22(\cpu|cpu|A_st_data[22]~q ),
	.A_mem_byte_en_2(\cpu|cpu|A_mem_byte_en[2]~q ),
	.A_st_data_23(\cpu|cpu|A_st_data[23]~q ),
	.A_st_data_24(\cpu|cpu|A_st_data[24]~q ),
	.A_mem_byte_en_3(\cpu|cpu|A_mem_byte_en[3]~q ),
	.A_st_data_25(\cpu|cpu|A_st_data[25]~q ),
	.A_st_data_31(\cpu|cpu|A_st_data[31]~q ),
	.A_st_data_21(\cpu|cpu|A_st_data[21]~q ),
	.A_st_data_11(\cpu|cpu|A_st_data[11]~q ),
	.A_mem_byte_en_1(\cpu|cpu|A_mem_byte_en[1]~q ),
	.A_st_data_28(\cpu|cpu|A_st_data[28]~q ),
	.A_st_data_10(\cpu|cpu|A_st_data[10]~q ),
	.A_st_data_27(\cpu|cpu|A_st_data[27]~q ),
	.A_st_data_8(\cpu|cpu|A_st_data[8]~q ),
	.A_st_data_9(\cpu|cpu|A_st_data[9]~q ),
	.A_st_data_26(\cpu|cpu|A_st_data[26]~q ),
	.A_st_data_20(\cpu|cpu|A_st_data[20]~q ),
	.A_st_data_19(\cpu|cpu|A_st_data[19]~q ),
	.A_st_data_17(\cpu|cpu|A_st_data[17]~q ),
	.A_st_data_30(\cpu|cpu|A_st_data[30]~q ),
	.A_st_data_18(\cpu|cpu|A_st_data[18]~q ),
	.A_st_data_15(\cpu|cpu|A_st_data[15]~q ),
	.A_st_data_12(\cpu|cpu|A_st_data[12]~q ),
	.A_st_data_13(\cpu|cpu|A_st_data[13]~q ),
	.A_st_data_14(\cpu|cpu|A_st_data[14]~q ),
	.A_st_data_29(\cpu|cpu|A_st_data[29]~q ),
	.src_data_26(\mm_interconnect_0|rsp_mux_001|src_data[26]~combout ),
	.src_data_25(\mm_interconnect_0|rsp_mux_001|src_data[25]~combout ),
	.src_data_24(\mm_interconnect_0|rsp_mux_001|src_data[24]~combout ),
	.src_data_23(\mm_interconnect_0|rsp_mux_001|src_data[23]~combout ),
	.src_data_22(\mm_interconnect_0|rsp_mux_001|src_data[22]~combout ),
	.src_data_11(\mm_interconnect_0|rsp_mux_001|src_data[1]~combout ),
	.src_data_01(\mm_interconnect_0|rsp_mux_001|src_data[0]~combout ),
	.src_data_21(\mm_interconnect_0|rsp_mux_001|src_data[2]~combout ),
	.src_data_31(\mm_interconnect_0|rsp_mux_001|src_data[3]~combout ),
	.src_data_4(\mm_interconnect_0|rsp_mux_001|src_data[4]~combout ),
	.src_data_5(\mm_interconnect_0|rsp_mux_001|src_data[5]~combout ),
	.src_data_28(\mm_interconnect_0|rsp_mux_001|src_data[28]~combout ),
	.src_data_311(\mm_interconnect_0|rsp_mux_001|src_data[31]~combout ),
	.src_data_27(\mm_interconnect_0|rsp_mux_001|src_data[27]~combout ),
	.src_data_29(\mm_interconnect_0|rsp_mux_001|src_data[29]~combout ),
	.src_data_30(\mm_interconnect_0|rsp_mux_001|src_data[30]~combout ),
	.src_data_111(\mm_interconnect_0|rsp_mux_001|src_data[11]~combout ),
	.src_data_12(\mm_interconnect_0|rsp_mux_001|src_data[12]~combout ),
	.src_data_13(\mm_interconnect_0|rsp_mux_001|src_data[13]~combout ),
	.src_data_14(\mm_interconnect_0|rsp_mux_001|src_data[14]~combout ),
	.src_data_15(\mm_interconnect_0|rsp_mux_001|src_data[15]~combout ),
	.src_data_16(\mm_interconnect_0|rsp_mux_001|src_data[16]~combout ),
	.src_payload46(\mm_interconnect_0|cmd_mux_002|src_payload~5_combout ),
	.src_data_9(\mm_interconnect_0|rsp_mux_001|src_data[9]~combout ),
	.src_data_211(\mm_interconnect_0|rsp_mux_001|src_data[21]~combout ),
	.src_data_6(\mm_interconnect_0|rsp_mux_001|src_data[6]~combout ),
	.src_data_8(\mm_interconnect_0|rsp_mux_001|src_data[8]~combout ),
	.src_data_17(\mm_interconnect_0|rsp_mux_001|src_data[17]~combout ),
	.src_data_18(\mm_interconnect_0|rsp_mux_001|src_data[18]~combout ),
	.src_data_10(\mm_interconnect_0|rsp_mux_001|src_data[10]~combout ),
	.src_data_7(\mm_interconnect_0|rsp_mux_001|src_data[7]~combout ),
	.src_data_20(\mm_interconnect_0|rsp_mux_001|src_data[20]~combout ),
	.src_data_19(\mm_interconnect_0|rsp_mux_001|src_data[19]~combout ),
	.src_payload47(\mm_interconnect_0|cmd_mux_002|src_payload~6_combout ),
	.src_data_34(\mm_interconnect_0|cmd_mux_002|src_data[34]~combout ),
	.src_payload48(\mm_interconnect_0|cmd_mux_002|src_payload~7_combout ),
	.src_payload49(\mm_interconnect_0|cmd_mux_002|src_payload~8_combout ),
	.src_payload50(\mm_interconnect_0|cmd_mux_002|src_payload~9_combout ),
	.src_payload51(\mm_interconnect_0|cmd_mux_002|src_payload~10_combout ),
	.src_payload52(\mm_interconnect_0|cmd_mux_002|src_payload~11_combout ),
	.src_payload53(\mm_interconnect_0|cmd_mux_002|src_payload~12_combout ),
	.src_payload54(\mm_interconnect_0|cmd_mux_002|src_payload~13_combout ),
	.src_payload55(\mm_interconnect_0|cmd_mux_002|src_payload~14_combout ),
	.src_payload56(\mm_interconnect_0|cmd_mux_002|src_payload~15_combout ),
	.src_data_35(\mm_interconnect_0|cmd_mux_002|src_data[35]~combout ),
	.src_payload57(\mm_interconnect_0|cmd_mux_002|src_payload~16_combout ),
	.src_payload58(\mm_interconnect_0|cmd_mux_002|src_payload~17_combout ),
	.src_payload59(\mm_interconnect_0|cmd_mux_002|src_payload~18_combout ),
	.src_payload60(\mm_interconnect_0|cmd_mux_002|src_payload~19_combout ),
	.src_payload61(\mm_interconnect_0|cmd_mux_002|src_payload~20_combout ),
	.src_payload62(\mm_interconnect_0|cmd_mux_002|src_payload~21_combout ),
	.src_payload63(\mm_interconnect_0|cmd_mux_002|src_payload~22_combout ),
	.src_data_33(\mm_interconnect_0|cmd_mux_002|src_data[33]~combout ),
	.src_payload64(\mm_interconnect_0|cmd_mux_002|src_payload~23_combout ),
	.src_payload65(\mm_interconnect_0|cmd_mux_002|src_payload~24_combout ),
	.src_payload66(\mm_interconnect_0|cmd_mux_002|src_payload~25_combout ),
	.src_payload67(\mm_interconnect_0|cmd_mux_002|src_payload~26_combout ),
	.src_payload68(\mm_interconnect_0|cmd_mux_002|src_payload~27_combout ),
	.src_payload69(\mm_interconnect_0|cmd_mux_002|src_payload~28_combout ),
	.src_payload70(\mm_interconnect_0|cmd_mux_002|src_payload~29_combout ),
	.src_payload71(\mm_interconnect_0|cmd_mux_002|src_payload~30_combout ),
	.src_payload72(\mm_interconnect_0|cmd_mux_002|src_payload~31_combout ),
	.src_payload73(\mm_interconnect_0|cmd_mux_002|src_payload~32_combout ),
	.altera_internal_jtag(\altera_internal_jtag~TCKUTAP ),
	.altera_internal_jtag1(\altera_internal_jtag~TDIUTAP ),
	.state_1(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.state_4(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.virtual_ir_scan_reg(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.state_3(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.state_8(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.splitter_nodes_receive_1_3(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_1[3]~q ),
	.irf_reg_0_2(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~q ),
	.irf_reg_1_2(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][1]~q ),
	.clk_clk(\clk_clk~input_o ));

first_nios2_system_first_nios2_system_camState1_1 camstate2(
	.readdata_0(\camstate2|readdata[0]~q ),
	.readdata_1(\camstate2|readdata[1]~q ),
	.readdata_2(\camstate2|readdata[2]~q ),
	.readdata_3(\camstate2|readdata[3]~q ),
	.readdata_4(\camstate2|readdata[4]~q ),
	.readdata_5(\camstate2|readdata[5]~q ),
	.Equal0(\camdata1|Equal0~0_combout ),
	.r_sync_rst(\rst_controller|r_sync_rst~q ),
	.clk_clk(\clk_clk~input_o ),
	.camstate2_external_connection_export_0(\camstate2_external_connection_export[0]~input_o ),
	.camstate2_external_connection_export_1(\camstate2_external_connection_export[1]~input_o ),
	.camstate2_external_connection_export_2(\camstate2_external_connection_export[2]~input_o ),
	.camstate2_external_connection_export_3(\camstate2_external_connection_export[3]~input_o ),
	.camstate2_external_connection_export_4(\camstate2_external_connection_export[4]~input_o ),
	.camstate2_external_connection_export_5(\camstate2_external_connection_export[5]~input_o ));

first_nios2_system_first_nios2_system_camState1 camstate1(
	.readdata_0(\camstate1|readdata[0]~q ),
	.readdata_1(\camstate1|readdata[1]~q ),
	.readdata_2(\camstate1|readdata[2]~q ),
	.readdata_3(\camstate1|readdata[3]~q ),
	.readdata_4(\camstate1|readdata[4]~q ),
	.readdata_5(\camstate1|readdata[5]~q ),
	.Equal0(\camdata1|Equal0~0_combout ),
	.r_sync_rst(\rst_controller|r_sync_rst~q ),
	.clk_clk(\clk_clk~input_o ),
	.camstate1_external_connection_export_0(\camstate1_external_connection_export[0]~input_o ),
	.camstate1_external_connection_export_1(\camstate1_external_connection_export[1]~input_o ),
	.camstate1_external_connection_export_2(\camstate1_external_connection_export[2]~input_o ),
	.camstate1_external_connection_export_3(\camstate1_external_connection_export[3]~input_o ),
	.camstate1_external_connection_export_4(\camstate1_external_connection_export[4]~input_o ),
	.camstate1_external_connection_export_5(\camstate1_external_connection_export[5]~input_o ));

first_nios2_system_first_nios2_system_camData1_1 camdata2(
	.readdata_0(\camdata2|readdata[0]~q ),
	.readdata_1(\camdata2|readdata[1]~q ),
	.readdata_2(\camdata2|readdata[2]~q ),
	.readdata_3(\camdata2|readdata[3]~q ),
	.readdata_4(\camdata2|readdata[4]~q ),
	.readdata_5(\camdata2|readdata[5]~q ),
	.readdata_6(\camdata2|readdata[6]~q ),
	.Equal0(\camdata1|Equal0~0_combout ),
	.r_sync_rst(\rst_controller|r_sync_rst~q ),
	.clk_clk(\clk_clk~input_o ),
	.camdata2_external_connection_export_0(\camdata2_external_connection_export[0]~input_o ),
	.camdata2_external_connection_export_1(\camdata2_external_connection_export[1]~input_o ),
	.camdata2_external_connection_export_2(\camdata2_external_connection_export[2]~input_o ),
	.camdata2_external_connection_export_3(\camdata2_external_connection_export[3]~input_o ),
	.camdata2_external_connection_export_4(\camdata2_external_connection_export[4]~input_o ),
	.camdata2_external_connection_export_5(\camdata2_external_connection_export[5]~input_o ),
	.camdata2_external_connection_export_6(\camdata2_external_connection_export[6]~input_o ));

first_nios2_system_first_nios2_system_camData1 camdata1(
	.readdata_0(\camdata1|readdata[0]~q ),
	.readdata_1(\camdata1|readdata[1]~q ),
	.readdata_2(\camdata1|readdata[2]~q ),
	.readdata_3(\camdata1|readdata[3]~q ),
	.readdata_4(\camdata1|readdata[4]~q ),
	.readdata_5(\camdata1|readdata[5]~q ),
	.readdata_6(\camdata1|readdata[6]~q ),
	.A_mem_baddr_3(\cpu|cpu|A_mem_baddr[3]~q ),
	.A_mem_baddr_2(\cpu|cpu|A_mem_baddr[2]~q ),
	.Equal0(\camdata1|Equal0~0_combout ),
	.r_sync_rst(\rst_controller|r_sync_rst~q ),
	.clk_clk(\clk_clk~input_o ),
	.camdata1_external_connection_export_0(\camdata1_external_connection_export[0]~input_o ),
	.camdata1_external_connection_export_1(\camdata1_external_connection_export[1]~input_o ),
	.camdata1_external_connection_export_2(\camdata1_external_connection_export[2]~input_o ),
	.camdata1_external_connection_export_3(\camdata1_external_connection_export[3]~input_o ),
	.camdata1_external_connection_export_4(\camdata1_external_connection_export[4]~input_o ),
	.camdata1_external_connection_export_5(\camdata1_external_connection_export[5]~input_o ),
	.camdata1_external_connection_export_6(\camdata1_external_connection_export[6]~input_o ));

first_nios2_system_first_nios2_system_sys_clk_timer sys_clk_timer(
	.writedata({\cpu|cpu|A_st_data[15]~q ,\cpu|cpu|A_st_data[14]~q ,\cpu|cpu|A_st_data[13]~q ,\cpu|cpu|A_st_data[12]~q ,\cpu|cpu|A_st_data[11]~q ,\cpu|cpu|A_st_data[10]~q ,\cpu|cpu|A_st_data[9]~q ,\cpu|cpu|A_st_data[8]~q ,\cpu|cpu|A_st_data[7]~q ,\cpu|cpu|A_st_data[6]~q ,
\cpu|cpu|A_st_data[5]~q ,\cpu|cpu|A_st_data[4]~q ,\cpu|cpu|A_st_data[3]~q ,\cpu|cpu|A_st_data[2]~q ,\cpu|cpu|A_st_data[1]~q ,\cpu|cpu|A_st_data[0]~q }),
	.A_mem_baddr_4(\cpu|cpu|A_mem_baddr[4]~q ),
	.clr_break_line(\cpu|cpu|clr_break_line~q ),
	.d_write(\cpu|cpu|d_write~q ),
	.A_mem_baddr_3(\cpu|cpu|A_mem_baddr[3]~q ),
	.A_mem_baddr_2(\cpu|cpu|A_mem_baddr[2]~q ),
	.reset_n(\rst_controller|r_sync_rst~q ),
	.Equal2(\mm_interconnect_0|router|Equal2~2_combout ),
	.wait_latency_counter_0(\mm_interconnect_0|sys_clk_timer_s1_translator|wait_latency_counter[0]~q ),
	.mem_used_1(\mm_interconnect_0|sys_clk_timer_s1_agent_rsp_fifo|mem_used[1]~q ),
	.wait_latency_counter_1(\mm_interconnect_0|sys_clk_timer_s1_translator|wait_latency_counter[1]~q ),
	.timeout_occurred1(\sys_clk_timer|timeout_occurred~q ),
	.control_register_0(\sys_clk_timer|control_register[0]~q ),
	.readdata_0(\sys_clk_timer|readdata[0]~q ),
	.readdata_1(\sys_clk_timer|readdata[1]~q ),
	.readdata_2(\sys_clk_timer|readdata[2]~q ),
	.readdata_3(\sys_clk_timer|readdata[3]~q ),
	.readdata_4(\sys_clk_timer|readdata[4]~q ),
	.readdata_5(\sys_clk_timer|readdata[5]~q ),
	.readdata_6(\sys_clk_timer|readdata[6]~q ),
	.readdata_7(\sys_clk_timer|readdata[7]~q ),
	.readdata_11(\sys_clk_timer|readdata[11]~q ),
	.readdata_10(\sys_clk_timer|readdata[10]~q ),
	.readdata_8(\sys_clk_timer|readdata[8]~q ),
	.readdata_9(\sys_clk_timer|readdata[9]~q ),
	.readdata_15(\sys_clk_timer|readdata[15]~q ),
	.readdata_12(\sys_clk_timer|readdata[12]~q ),
	.readdata_13(\sys_clk_timer|readdata[13]~q ),
	.readdata_14(\sys_clk_timer|readdata[14]~q ),
	.clk(\clk_clk~input_o ));

first_nios2_system_first_nios2_system_download1_2 start(
	.data_out1(\start|data_out~q ),
	.A_st_data_0(\cpu|cpu|A_st_data[0]~q ),
	.clr_break_line(\cpu|cpu|clr_break_line~q ),
	.d_write(\cpu|cpu|d_write~q ),
	.Equal0(\camdata1|Equal0~0_combout ),
	.reset_n(\rst_controller|r_sync_rst~q ),
	.wait_latency_counter_1(\mm_interconnect_0|start_s1_translator|wait_latency_counter[1]~q ),
	.m0_write(\mm_interconnect_0|start_s1_agent|m0_write~0_combout ),
	.wait_latency_counter_0(\mm_interconnect_0|start_s1_translator|wait_latency_counter[0]~q ),
	.clk(\clk_clk~input_o ));

first_nios2_system_first_nios2_system_rtd1_1 rtd2(
	.readdata_0(\rtd2|readdata[0]~q ),
	.Equal0(\camdata1|Equal0~0_combout ),
	.r_sync_rst(\rst_controller|r_sync_rst~q ),
	.clk_clk(\clk_clk~input_o ),
	.rtd2_external_connection_export(\rtd2_external_connection_export~input_o ));

first_nios2_system_first_nios2_system_rtd1 rtd1(
	.readdata_0(\rtd1|readdata[0]~q ),
	.Equal0(\camdata1|Equal0~0_combout ),
	.r_sync_rst(\rst_controller|r_sync_rst~q ),
	.clk_clk(\clk_clk~input_o ),
	.rtd1_external_connection_export(\rtd1_external_connection_export~input_o ));

first_nios2_system_first_nios2_system_onchip_mem onchip_mem(
	.q_a_0(\onchip_mem|the_altsyncram|auto_generated|q_a[0] ),
	.q_a_1(\onchip_mem|the_altsyncram|auto_generated|q_a[1] ),
	.q_a_2(\onchip_mem|the_altsyncram|auto_generated|q_a[2] ),
	.q_a_3(\onchip_mem|the_altsyncram|auto_generated|q_a[3] ),
	.q_a_4(\onchip_mem|the_altsyncram|auto_generated|q_a[4] ),
	.q_a_5(\onchip_mem|the_altsyncram|auto_generated|q_a[5] ),
	.q_a_6(\onchip_mem|the_altsyncram|auto_generated|q_a[6] ),
	.q_a_7(\onchip_mem|the_altsyncram|auto_generated|q_a[7] ),
	.q_a_22(\onchip_mem|the_altsyncram|auto_generated|q_a[22] ),
	.q_a_23(\onchip_mem|the_altsyncram|auto_generated|q_a[23] ),
	.q_a_24(\onchip_mem|the_altsyncram|auto_generated|q_a[24] ),
	.q_a_25(\onchip_mem|the_altsyncram|auto_generated|q_a[25] ),
	.q_a_31(\onchip_mem|the_altsyncram|auto_generated|q_a[31] ),
	.q_a_21(\onchip_mem|the_altsyncram|auto_generated|q_a[21] ),
	.q_a_11(\onchip_mem|the_altsyncram|auto_generated|q_a[11] ),
	.q_a_28(\onchip_mem|the_altsyncram|auto_generated|q_a[28] ),
	.q_a_10(\onchip_mem|the_altsyncram|auto_generated|q_a[10] ),
	.q_a_27(\onchip_mem|the_altsyncram|auto_generated|q_a[27] ),
	.q_a_8(\onchip_mem|the_altsyncram|auto_generated|q_a[8] ),
	.q_a_9(\onchip_mem|the_altsyncram|auto_generated|q_a[9] ),
	.q_a_26(\onchip_mem|the_altsyncram|auto_generated|q_a[26] ),
	.q_a_20(\onchip_mem|the_altsyncram|auto_generated|q_a[20] ),
	.q_a_19(\onchip_mem|the_altsyncram|auto_generated|q_a[19] ),
	.q_a_17(\onchip_mem|the_altsyncram|auto_generated|q_a[17] ),
	.q_a_30(\onchip_mem|the_altsyncram|auto_generated|q_a[30] ),
	.q_a_18(\onchip_mem|the_altsyncram|auto_generated|q_a[18] ),
	.q_a_16(\onchip_mem|the_altsyncram|auto_generated|q_a[16] ),
	.q_a_15(\onchip_mem|the_altsyncram|auto_generated|q_a[15] ),
	.q_a_12(\onchip_mem|the_altsyncram|auto_generated|q_a[12] ),
	.q_a_13(\onchip_mem|the_altsyncram|auto_generated|q_a[13] ),
	.q_a_14(\onchip_mem|the_altsyncram|auto_generated|q_a[14] ),
	.q_a_29(\onchip_mem|the_altsyncram|auto_generated|q_a[29] ),
	.d_write(\cpu|cpu|d_write~q ),
	.mem_used_1(\mm_interconnect_0|onchip_mem_s1_agent_rsp_fifo|mem_used[1]~q ),
	.saved_grant_0(\mm_interconnect_0|cmd_mux_003|saved_grant[0]~q ),
	.WideOr1(\mm_interconnect_0|cmd_mux_003|WideOr1~combout ),
	.r_early_rst(\rst_controller|r_early_rst~q ),
	.src_payload(\mm_interconnect_0|cmd_mux_003|src_payload~0_combout ),
	.src_data_38(\mm_interconnect_0|cmd_mux_003|src_data[38]~combout ),
	.src_data_39(\mm_interconnect_0|cmd_mux_003|src_data[39]~combout ),
	.src_data_40(\mm_interconnect_0|cmd_mux_003|src_data[40]~combout ),
	.src_data_41(\mm_interconnect_0|cmd_mux_003|src_data[41]~combout ),
	.src_data_42(\mm_interconnect_0|cmd_mux_003|src_data[42]~combout ),
	.src_data_43(\mm_interconnect_0|cmd_mux_003|src_data[43]~combout ),
	.src_data_44(\mm_interconnect_0|cmd_mux_003|src_data[44]~combout ),
	.src_data_45(\mm_interconnect_0|cmd_mux_003|src_data[45]~combout ),
	.src_data_46(\mm_interconnect_0|cmd_mux_003|src_data[46]~combout ),
	.src_data_47(\mm_interconnect_0|cmd_mux_003|src_data[47]~combout ),
	.src_data_48(\mm_interconnect_0|cmd_mux_003|src_data[48]~combout ),
	.src_data_49(\mm_interconnect_0|cmd_mux_003|src_data[49]~combout ),
	.src_data_50(\mm_interconnect_0|cmd_mux_003|src_data[50]~combout ),
	.src_data_32(\mm_interconnect_0|cmd_mux_003|src_data[32]~combout ),
	.src_payload1(\mm_interconnect_0|cmd_mux_003|src_payload~1_combout ),
	.src_payload2(\mm_interconnect_0|cmd_mux_003|src_payload~2_combout ),
	.src_payload3(\mm_interconnect_0|cmd_mux_003|src_payload~3_combout ),
	.src_payload4(\mm_interconnect_0|cmd_mux_003|src_payload~4_combout ),
	.src_payload5(\mm_interconnect_0|cmd_mux_003|src_payload~5_combout ),
	.src_payload6(\mm_interconnect_0|cmd_mux_003|src_payload~6_combout ),
	.src_payload7(\mm_interconnect_0|cmd_mux_003|src_payload~7_combout ),
	.src_payload8(\mm_interconnect_0|cmd_mux_003|src_payload~8_combout ),
	.src_data_34(\mm_interconnect_0|cmd_mux_003|src_data[34]~combout ),
	.src_payload9(\mm_interconnect_0|cmd_mux_003|src_payload~9_combout ),
	.src_payload10(\mm_interconnect_0|cmd_mux_003|src_payload~10_combout ),
	.src_data_35(\mm_interconnect_0|cmd_mux_003|src_data[35]~combout ),
	.src_payload11(\mm_interconnect_0|cmd_mux_003|src_payload~11_combout ),
	.src_payload12(\mm_interconnect_0|cmd_mux_003|src_payload~12_combout ),
	.src_payload13(\mm_interconnect_0|cmd_mux_003|src_payload~13_combout ),
	.src_payload14(\mm_interconnect_0|cmd_mux_003|src_payload~14_combout ),
	.src_data_33(\mm_interconnect_0|cmd_mux_003|src_data[33]~combout ),
	.src_payload15(\mm_interconnect_0|cmd_mux_003|src_payload~15_combout ),
	.src_payload16(\mm_interconnect_0|cmd_mux_003|src_payload~16_combout ),
	.src_payload17(\mm_interconnect_0|cmd_mux_003|src_payload~17_combout ),
	.src_payload18(\mm_interconnect_0|cmd_mux_003|src_payload~18_combout ),
	.src_payload19(\mm_interconnect_0|cmd_mux_003|src_payload~19_combout ),
	.src_payload20(\mm_interconnect_0|cmd_mux_003|src_payload~20_combout ),
	.src_payload21(\mm_interconnect_0|cmd_mux_003|src_payload~21_combout ),
	.src_payload22(\mm_interconnect_0|cmd_mux_003|src_payload~22_combout ),
	.src_payload23(\mm_interconnect_0|cmd_mux_003|src_payload~23_combout ),
	.src_payload24(\mm_interconnect_0|cmd_mux_003|src_payload~24_combout ),
	.src_payload25(\mm_interconnect_0|cmd_mux_003|src_payload~25_combout ),
	.src_payload26(\mm_interconnect_0|cmd_mux_003|src_payload~26_combout ),
	.src_payload27(\mm_interconnect_0|cmd_mux_003|src_payload~27_combout ),
	.src_payload28(\mm_interconnect_0|cmd_mux_003|src_payload~28_combout ),
	.src_payload29(\mm_interconnect_0|cmd_mux_003|src_payload~29_combout ),
	.src_payload30(\mm_interconnect_0|cmd_mux_003|src_payload~30_combout ),
	.src_payload31(\mm_interconnect_0|cmd_mux_003|src_payload~31_combout ),
	.clk_clk(\clk_clk~input_o ));

first_nios2_system_first_nios2_system_leds leds(
	.data_out_0(\leds|data_out[0]~q ),
	.data_out_1(\leds|data_out[1]~q ),
	.data_out_2(\leds|data_out[2]~q ),
	.data_out_3(\leds|data_out[3]~q ),
	.data_out_4(\leds|data_out[4]~q ),
	.data_out_5(\leds|data_out[5]~q ),
	.data_out_6(\leds|data_out[6]~q ),
	.data_out_7(\leds|data_out[7]~q ),
	.writedata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\cpu|cpu|A_st_data[7]~q ,\cpu|cpu|A_st_data[6]~q ,\cpu|cpu|A_st_data[5]~q ,\cpu|cpu|A_st_data[4]~q ,\cpu|cpu|A_st_data[3]~q ,\cpu|cpu|A_st_data[2]~q ,\cpu|cpu|A_st_data[1]~q ,
\cpu|cpu|A_st_data[0]~q }),
	.clr_break_line(\cpu|cpu|clr_break_line~q ),
	.d_write(\cpu|cpu|d_write~q ),
	.Equal0(\camdata1|Equal0~0_combout ),
	.reset_n(\rst_controller|r_sync_rst~q ),
	.wait_latency_counter_1(\mm_interconnect_0|leds_s1_translator|wait_latency_counter[1]~q ),
	.mem_used_1(\mm_interconnect_0|leds_s1_agent_rsp_fifo|mem_used[1]~q ),
	.Equal16(\mm_interconnect_0|router|Equal16~0_combout ),
	.wait_latency_counter_0(\mm_interconnect_0|leds_s1_translator|wait_latency_counter[0]~q ),
	.clk(\clk_clk~input_o ));

first_nios2_system_first_nios2_system_jtag_uart jtag_uart(
	.q_b_0(\jtag_uart|the_first_nios2_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[0] ),
	.q_b_1(\jtag_uart|the_first_nios2_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[1] ),
	.q_b_2(\jtag_uart|the_first_nios2_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[2] ),
	.q_b_3(\jtag_uart|the_first_nios2_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[3] ),
	.q_b_4(\jtag_uart|the_first_nios2_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[4] ),
	.q_b_5(\jtag_uart|the_first_nios2_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.q_b_6(\jtag_uart|the_first_nios2_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.q_b_7(\jtag_uart|the_first_nios2_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.Add1(\jtag_uart|Add1~1_sumout ),
	.Add11(\jtag_uart|Add1~5_sumout ),
	.Add12(\jtag_uart|Add1~9_sumout ),
	.Add13(\jtag_uart|Add1~13_sumout ),
	.Add14(\jtag_uart|Add1~17_sumout ),
	.Add15(\jtag_uart|Add1~21_sumout ),
	.Add16(\jtag_uart|Add1~25_sumout ),
	.tdo(\jtag_uart|first_nios2_system_jtag_uart_alt_jtag_atlantic|tdo~q ),
	.A_st_data_0(\cpu|cpu|A_st_data[0]~q ),
	.A_mem_baddr_4(\cpu|cpu|A_mem_baddr[4]~q ),
	.Equal1(\mm_interconnect_0|router|Equal1~0_combout ),
	.Equal2(\mm_interconnect_0|router|Equal2~0_combout ),
	.clr_break_line(\cpu|cpu|clr_break_line~q ),
	.d_write(\cpu|cpu|d_write~q ),
	.A_mem_baddr_3(\cpu|cpu|A_mem_baddr[3]~q ),
	.A_mem_baddr_2(\cpu|cpu|A_mem_baddr[2]~q ),
	.r_sync_rst(\rst_controller|r_sync_rst~q ),
	.A_st_data_1(\cpu|cpu|A_st_data[1]~q ),
	.A_st_data_2(\cpu|cpu|A_st_data[2]~q ),
	.A_st_data_3(\cpu|cpu|A_st_data[3]~q ),
	.A_st_data_4(\cpu|cpu|A_st_data[4]~q ),
	.A_st_data_5(\cpu|cpu|A_st_data[5]~q ),
	.A_st_data_6(\cpu|cpu|A_st_data[6]~q ),
	.A_st_data_7(\cpu|cpu|A_st_data[7]~q ),
	.read_latency_shift_reg(\mm_interconnect_0|download1_s1_translator|read_latency_shift_reg~0_combout ),
	.cp_valid(\mm_interconnect_0|cpu_data_master_agent|cp_valid~0_combout ),
	.always1(\mm_interconnect_0|router|always1~2_combout ),
	.av_waitrequest1(\jtag_uart|av_waitrequest~q ),
	.mem_used_1(\mm_interconnect_0|jtag_uart_avalon_jtag_slave_agent_rsp_fifo|mem_used[1]~q ),
	.av_waitrequest2(\jtag_uart|av_waitrequest~0_combout ),
	.ien_AE1(\jtag_uart|ien_AE~q ),
	.av_readdata_9(\jtag_uart|av_readdata[9]~combout ),
	.ien_AF1(\jtag_uart|ien_AF~q ),
	.av_readdata_8(\jtag_uart|av_readdata[8]~0_combout ),
	.b_full(\jtag_uart|the_first_nios2_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|b_full~q ),
	.b_full1(\jtag_uart|the_first_nios2_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|b_full~q ),
	.b_non_empty(\jtag_uart|the_first_nios2_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|b_non_empty~q ),
	.read_01(\jtag_uart|read_0~q ),
	.counter_reg_bit_0(\jtag_uart|the_first_nios2_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\jtag_uart|the_first_nios2_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[1]~q ),
	.counter_reg_bit_4(\jtag_uart|the_first_nios2_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[4]~q ),
	.counter_reg_bit_3(\jtag_uart|the_first_nios2_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[3]~q ),
	.counter_reg_bit_2(\jtag_uart|the_first_nios2_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[2]~q ),
	.counter_reg_bit_5(\jtag_uart|the_first_nios2_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[5]~q ),
	.A_st_data_10(\cpu|cpu|A_st_data[10]~q ),
	.ac1(\jtag_uart|ac~q ),
	.rvalid1(\jtag_uart|rvalid~q ),
	.woverflow1(\jtag_uart|woverflow~q ),
	.altera_internal_jtag(\altera_internal_jtag~TCKUTAP ),
	.altera_internal_jtag1(\altera_internal_jtag~TDIUTAP ),
	.state_4(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.splitter_nodes_receive_0_3(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ),
	.virtual_ir_scan_reg(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.clr_reg(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.state_3(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.state_8(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.irf_reg_0_1(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.clk_clk(\clk_clk~input_o ));

first_nios2_system_first_nios2_system_hex1_1 hex2(
	.data_out_0(\hex2|data_out[0]~q ),
	.data_out_1(\hex2|data_out[1]~q ),
	.data_out_2(\hex2|data_out[2]~q ),
	.data_out_3(\hex2|data_out[3]~q ),
	.data_out_4(\hex2|data_out[4]~q ),
	.data_out_5(\hex2|data_out[5]~q ),
	.data_out_6(\hex2|data_out[6]~q ),
	.writedata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\cpu|cpu|A_st_data[6]~q ,\cpu|cpu|A_st_data[5]~q ,\cpu|cpu|A_st_data[4]~q ,\cpu|cpu|A_st_data[3]~q ,\cpu|cpu|A_st_data[2]~q ,\cpu|cpu|A_st_data[1]~q ,\cpu|cpu|A_st_data[0]~q }),
	.A_mem_baddr_7(\cpu|cpu|A_mem_baddr[7]~q ),
	.clr_break_line(\cpu|cpu|clr_break_line~q ),
	.d_write(\cpu|cpu|d_write~q ),
	.Equal0(\camdata1|Equal0~0_combout ),
	.reset_n(\rst_controller|r_sync_rst~q ),
	.wait_latency_counter_1(\mm_interconnect_0|hex2_s1_translator|wait_latency_counter[1]~q ),
	.mem_used_1(\mm_interconnect_0|hex2_s1_agent_rsp_fifo|mem_used[1]~q ),
	.always1(\mm_interconnect_0|router|always1~0_combout ),
	.wait_latency_counter_0(\mm_interconnect_0|hex2_s1_translator|wait_latency_counter[0]~q ),
	.clk(\clk_clk~input_o ));

first_nios2_system_first_nios2_system_hex1 hex1(
	.data_out_0(\hex1|data_out[0]~q ),
	.data_out_1(\hex1|data_out[1]~q ),
	.data_out_2(\hex1|data_out[2]~q ),
	.data_out_3(\hex1|data_out[3]~q ),
	.data_out_4(\hex1|data_out[4]~q ),
	.data_out_5(\hex1|data_out[5]~q ),
	.data_out_6(\hex1|data_out[6]~q ),
	.writedata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\cpu|cpu|A_st_data[6]~q ,\cpu|cpu|A_st_data[5]~q ,\cpu|cpu|A_st_data[4]~q ,\cpu|cpu|A_st_data[3]~q ,\cpu|cpu|A_st_data[2]~q ,\cpu|cpu|A_st_data[1]~q ,\cpu|cpu|A_st_data[0]~q }),
	.clr_break_line(\cpu|cpu|clr_break_line~q ),
	.d_write(\cpu|cpu|d_write~q ),
	.Equal0(\camdata1|Equal0~0_combout ),
	.reset_n(\rst_controller|r_sync_rst~q ),
	.wait_latency_counter_1(\mm_interconnect_0|hex1_s1_translator|wait_latency_counter[1]~q ),
	.mem_used_1(\mm_interconnect_0|hex1_s1_agent_rsp_fifo|mem_used[1]~q ),
	.Equal6(\mm_interconnect_0|router|Equal6~1_combout ),
	.wait_latency_counter_0(\mm_interconnect_0|hex1_s1_translator|wait_latency_counter[0]~q ),
	.clk(\clk_clk~input_o ));

first_nios2_system_first_nios2_system_download1_1 download2(
	.data_out1(\download2|data_out~q ),
	.A_st_data_0(\cpu|cpu|A_st_data[0]~q ),
	.clr_break_line(\cpu|cpu|clr_break_line~q ),
	.d_write(\cpu|cpu|d_write~q ),
	.Equal0(\camdata1|Equal0~0_combout ),
	.reset_n(\rst_controller|r_sync_rst~q ),
	.write(\mm_interconnect_0|download2_s1_agent_rsp_fifo|write~0_combout ),
	.wait_latency_counter_0(\mm_interconnect_0|download2_s1_translator|wait_latency_counter[0]~q ),
	.clk(\clk_clk~input_o ));

first_nios2_system_first_nios2_system_download1 download1(
	.data_out1(\download1|data_out~q ),
	.A_st_data_0(\cpu|cpu|A_st_data[0]~q ),
	.mem_used_1(\mm_interconnect_0|download1_s1_agent_rsp_fifo|mem_used[1]~q ),
	.Equal15(\mm_interconnect_0|router|Equal15~1_combout ),
	.always0(\download1|always0~0_combout ),
	.clr_break_line(\cpu|cpu|clr_break_line~q ),
	.wait_latency_counter_1(\mm_interconnect_0|download1_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\mm_interconnect_0|download1_s1_translator|wait_latency_counter[0]~q ),
	.d_write(\cpu|cpu|d_write~q ),
	.Equal0(\camdata1|Equal0~0_combout ),
	.reset_n(\rst_controller|r_sync_rst~q ),
	.clk(\clk_clk~input_o ));

first_nios2_system_first_nios2_system_mm_interconnect_0 mm_interconnect_0(
	.q_a_0(\onchip_mem|the_altsyncram|auto_generated|q_a[0] ),
	.q_a_1(\onchip_mem|the_altsyncram|auto_generated|q_a[1] ),
	.q_a_2(\onchip_mem|the_altsyncram|auto_generated|q_a[2] ),
	.q_a_3(\onchip_mem|the_altsyncram|auto_generated|q_a[3] ),
	.q_a_4(\onchip_mem|the_altsyncram|auto_generated|q_a[4] ),
	.q_a_5(\onchip_mem|the_altsyncram|auto_generated|q_a[5] ),
	.q_a_6(\onchip_mem|the_altsyncram|auto_generated|q_a[6] ),
	.q_a_7(\onchip_mem|the_altsyncram|auto_generated|q_a[7] ),
	.av_readdata_pre_22(\mm_interconnect_0|jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[22]~q ),
	.q_a_22(\onchip_mem|the_altsyncram|auto_generated|q_a[22] ),
	.q_a_23(\onchip_mem|the_altsyncram|auto_generated|q_a[23] ),
	.q_a_24(\onchip_mem|the_altsyncram|auto_generated|q_a[24] ),
	.q_a_25(\onchip_mem|the_altsyncram|auto_generated|q_a[25] ),
	.q_a_31(\onchip_mem|the_altsyncram|auto_generated|q_a[31] ),
	.q_a_21(\onchip_mem|the_altsyncram|auto_generated|q_a[21] ),
	.q_a_11(\onchip_mem|the_altsyncram|auto_generated|q_a[11] ),
	.q_a_28(\onchip_mem|the_altsyncram|auto_generated|q_a[28] ),
	.q_a_10(\onchip_mem|the_altsyncram|auto_generated|q_a[10] ),
	.q_a_27(\onchip_mem|the_altsyncram|auto_generated|q_a[27] ),
	.q_a_8(\onchip_mem|the_altsyncram|auto_generated|q_a[8] ),
	.q_a_9(\onchip_mem|the_altsyncram|auto_generated|q_a[9] ),
	.q_a_26(\onchip_mem|the_altsyncram|auto_generated|q_a[26] ),
	.av_readdata_pre_20(\mm_interconnect_0|jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[20]~q ),
	.q_a_20(\onchip_mem|the_altsyncram|auto_generated|q_a[20] ),
	.av_readdata_pre_19(\mm_interconnect_0|jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[19]~q ),
	.q_a_19(\onchip_mem|the_altsyncram|auto_generated|q_a[19] ),
	.q_a_17(\onchip_mem|the_altsyncram|auto_generated|q_a[17] ),
	.q_a_30(\onchip_mem|the_altsyncram|auto_generated|q_a[30] ),
	.q_a_18(\onchip_mem|the_altsyncram|auto_generated|q_a[18] ),
	.q_a_16(\onchip_mem|the_altsyncram|auto_generated|q_a[16] ),
	.q_a_15(\onchip_mem|the_altsyncram|auto_generated|q_a[15] ),
	.q_a_12(\onchip_mem|the_altsyncram|auto_generated|q_a[12] ),
	.q_a_13(\onchip_mem|the_altsyncram|auto_generated|q_a[13] ),
	.q_a_14(\onchip_mem|the_altsyncram|auto_generated|q_a[14] ),
	.q_a_29(\onchip_mem|the_altsyncram|auto_generated|q_a[29] ),
	.readdata_0(\cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[0]~q ),
	.readdata_01(\camstate2|readdata[0]~q ),
	.readdata_02(\tenout1|readdata[0]~q ),
	.readdata_03(\tenout2|readdata[0]~q ),
	.readdata_04(\camstate1|readdata[0]~q ),
	.readdata_05(\rtd2|readdata[0]~q ),
	.readdata_06(\rtd1|readdata[0]~q ),
	.q_b_0(\jtag_uart|the_first_nios2_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[0] ),
	.readdata_07(\camdata1|readdata[0]~q ),
	.readdata_08(\camdata2|readdata[0]~q ),
	.readdata_1(\tenout2|readdata[1]~q ),
	.readdata_11(\cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[1]~q ),
	.readdata_12(\camdata1|readdata[1]~q ),
	.readdata_13(\camstate2|readdata[1]~q ),
	.q_b_1(\jtag_uart|the_first_nios2_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[1] ),
	.readdata_14(\camdata2|readdata[1]~q ),
	.readdata_15(\camstate1|readdata[1]~q ),
	.readdata_16(\tenout1|readdata[1]~q ),
	.readdata_2(\tenout2|readdata[2]~q ),
	.readdata_21(\cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[2]~q ),
	.readdata_22(\camdata1|readdata[2]~q ),
	.readdata_23(\camstate2|readdata[2]~q ),
	.q_b_2(\jtag_uart|the_first_nios2_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[2] ),
	.readdata_24(\camdata2|readdata[2]~q ),
	.readdata_25(\camstate1|readdata[2]~q ),
	.readdata_26(\tenout1|readdata[2]~q ),
	.readdata_3(\camdata2|readdata[3]~q ),
	.readdata_31(\tenout2|readdata[3]~q ),
	.readdata_32(\cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[3]~q ),
	.readdata_33(\camdata1|readdata[3]~q ),
	.readdata_34(\tenout1|readdata[3]~q ),
	.q_b_3(\jtag_uart|the_first_nios2_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[3] ),
	.readdata_35(\camstate1|readdata[3]~q ),
	.readdata_36(\camstate2|readdata[3]~q ),
	.q_b_4(\jtag_uart|the_first_nios2_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[4] ),
	.readdata_4(\cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[4]~q ),
	.readdata_41(\camdata1|readdata[4]~q ),
	.readdata_42(\camdata2|readdata[4]~q ),
	.readdata_43(\camstate1|readdata[4]~q ),
	.readdata_44(\camstate2|readdata[4]~q ),
	.readdata_5(\cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[5]~q ),
	.readdata_51(\camdata1|readdata[5]~q ),
	.readdata_52(\camdata2|readdata[5]~q ),
	.q_b_5(\jtag_uart|the_first_nios2_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.readdata_53(\camstate1|readdata[5]~q ),
	.readdata_54(\camstate2|readdata[5]~q ),
	.readdata_6(\camdata1|readdata[6]~q ),
	.q_b_6(\jtag_uart|the_first_nios2_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.readdata_61(\cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[6]~q ),
	.readdata_62(\camdata2|readdata[6]~q ),
	.q_b_7(\jtag_uart|the_first_nios2_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.readdata_7(\cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[7]~q ),
	.Add1(\jtag_uart|Add1~1_sumout ),
	.readdata_221(\cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[22]~q ),
	.readdata_231(\cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[23]~q ),
	.readdata_241(\cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[24]~q ),
	.readdata_251(\cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[25]~q ),
	.readdata_311(\cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[31]~q ),
	.readdata_211(\cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[21]~q ),
	.Add11(\jtag_uart|Add1~5_sumout ),
	.readdata_111(\cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[11]~q ),
	.readdata_28(\cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[28]~q ),
	.readdata_10(\cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[10]~q ),
	.readdata_27(\cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[27]~q ),
	.readdata_8(\cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[8]~q ),
	.readdata_9(\cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[9]~q ),
	.readdata_261(\cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[26]~q ),
	.Add12(\jtag_uart|Add1~9_sumout ),
	.readdata_20(\cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[20]~q ),
	.Add13(\jtag_uart|Add1~13_sumout ),
	.readdata_19(\cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[19]~q ),
	.readdata_17(\cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[17]~q ),
	.Add14(\jtag_uart|Add1~17_sumout ),
	.readdata_30(\cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[30]~q ),
	.readdata_18(\cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[18]~q ),
	.Add15(\jtag_uart|Add1~21_sumout ),
	.readdata_161(\cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[16]~q ),
	.Add16(\jtag_uart|Add1~25_sumout ),
	.readdata_151(\cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[15]~q ),
	.readdata_121(\cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[12]~q ),
	.readdata_131(\cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[13]~q ),
	.readdata_141(\cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[14]~q ),
	.readdata_29(\cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|readdata[29]~q ),
	.data_out(\download1|data_out~q ),
	.data_out1(\download2|data_out~q ),
	.data_out_0(\hex1|data_out[0]~q ),
	.data_out_1(\hex1|data_out[1]~q ),
	.data_out_2(\hex1|data_out[2]~q ),
	.data_out_3(\hex1|data_out[3]~q ),
	.data_out_4(\hex1|data_out[4]~q ),
	.data_out_5(\hex1|data_out[5]~q ),
	.data_out_6(\hex1|data_out[6]~q ),
	.data_out_01(\hex2|data_out[0]~q ),
	.data_out_11(\hex2|data_out[1]~q ),
	.data_out_21(\hex2|data_out[2]~q ),
	.data_out_31(\hex2|data_out[3]~q ),
	.data_out_41(\hex2|data_out[4]~q ),
	.data_out_51(\hex2|data_out[5]~q ),
	.data_out_61(\hex2|data_out[6]~q ),
	.data_out_02(\leds|data_out[0]~q ),
	.data_out_12(\leds|data_out[1]~q ),
	.data_out_22(\leds|data_out[2]~q ),
	.data_out_32(\leds|data_out[3]~q ),
	.data_out_42(\leds|data_out[4]~q ),
	.data_out_52(\leds|data_out[5]~q ),
	.data_out_62(\leds|data_out[6]~q ),
	.data_out_7(\leds|data_out[7]~q ),
	.data_out2(\start|data_out~q ),
	.A_st_data_0(\cpu|cpu|A_st_data[0]~q ),
	.mem_used_1(\mm_interconnect_0|download1_s1_agent_rsp_fifo|mem_used[1]~q ),
	.A_mem_baddr_4(\cpu|cpu|A_mem_baddr[4]~q ),
	.A_mem_baddr_5(\cpu|cpu|A_mem_baddr[5]~q ),
	.A_mem_baddr_8(\cpu|cpu|A_mem_baddr[8]~q ),
	.A_mem_baddr_16(\cpu|cpu|A_mem_baddr[16]~q ),
	.A_mem_baddr_15(\cpu|cpu|A_mem_baddr[15]~q ),
	.A_mem_baddr_14(\cpu|cpu|A_mem_baddr[14]~q ),
	.A_mem_baddr_13(\cpu|cpu|A_mem_baddr[13]~q ),
	.Equal1(\mm_interconnect_0|router|Equal1~0_combout ),
	.A_mem_baddr_12(\cpu|cpu|A_mem_baddr[12]~q ),
	.A_mem_baddr_11(\cpu|cpu|A_mem_baddr[11]~q ),
	.A_mem_baddr_10(\cpu|cpu|A_mem_baddr[10]~q ),
	.A_mem_baddr_9(\cpu|cpu|A_mem_baddr[9]~q ),
	.Equal2(\mm_interconnect_0|router|Equal2~0_combout ),
	.A_mem_baddr_7(\cpu|cpu|A_mem_baddr[7]~q ),
	.A_mem_baddr_6(\cpu|cpu|A_mem_baddr[6]~q ),
	.Equal15(\mm_interconnect_0|router|Equal15~1_combout ),
	.always0(\download1|always0~0_combout ),
	.clr_break_line(\cpu|cpu|clr_break_line~q ),
	.wait_latency_counter_1(\mm_interconnect_0|download1_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\mm_interconnect_0|download1_s1_translator|wait_latency_counter[0]~q ),
	.d_write(\cpu|cpu|d_write~q ),
	.A_mem_baddr_3(\cpu|cpu|A_mem_baddr[3]~q ),
	.A_mem_baddr_2(\cpu|cpu|A_mem_baddr[2]~q ),
	.Equal0(\camdata1|Equal0~0_combout ),
	.r_sync_rst(\rst_controller|r_sync_rst~q ),
	.write(\mm_interconnect_0|download2_s1_agent_rsp_fifo|write~0_combout ),
	.wait_latency_counter_01(\mm_interconnect_0|download2_s1_translator|wait_latency_counter[0]~q ),
	.wait_latency_counter_11(\mm_interconnect_0|hex1_s1_translator|wait_latency_counter[1]~q ),
	.mem_used_11(\mm_interconnect_0|hex1_s1_agent_rsp_fifo|mem_used[1]~q ),
	.Equal6(\mm_interconnect_0|router|Equal6~1_combout ),
	.wait_latency_counter_02(\mm_interconnect_0|hex1_s1_translator|wait_latency_counter[0]~q ),
	.A_st_data_1(\cpu|cpu|A_st_data[1]~q ),
	.A_st_data_2(\cpu|cpu|A_st_data[2]~q ),
	.A_st_data_3(\cpu|cpu|A_st_data[3]~q ),
	.A_st_data_4(\cpu|cpu|A_st_data[4]~q ),
	.A_st_data_5(\cpu|cpu|A_st_data[5]~q ),
	.A_st_data_6(\cpu|cpu|A_st_data[6]~q ),
	.wait_latency_counter_12(\mm_interconnect_0|hex2_s1_translator|wait_latency_counter[1]~q ),
	.mem_used_12(\mm_interconnect_0|hex2_s1_agent_rsp_fifo|mem_used[1]~q ),
	.always1(\mm_interconnect_0|router|always1~0_combout ),
	.wait_latency_counter_03(\mm_interconnect_0|hex2_s1_translator|wait_latency_counter[0]~q ),
	.wait_latency_counter_13(\mm_interconnect_0|leds_s1_translator|wait_latency_counter[1]~q ),
	.mem_used_13(\mm_interconnect_0|leds_s1_agent_rsp_fifo|mem_used[1]~q ),
	.Equal16(\mm_interconnect_0|router|Equal16~0_combout ),
	.wait_latency_counter_04(\mm_interconnect_0|leds_s1_translator|wait_latency_counter[0]~q ),
	.A_st_data_7(\cpu|cpu|A_st_data[7]~q ),
	.wait_latency_counter_14(\mm_interconnect_0|start_s1_translator|wait_latency_counter[1]~q ),
	.m0_write(\mm_interconnect_0|start_s1_agent|m0_write~0_combout ),
	.wait_latency_counter_05(\mm_interconnect_0|start_s1_translator|wait_latency_counter[0]~q ),
	.d_read(\cpu|cpu|d_read~q ),
	.read_latency_shift_reg(\mm_interconnect_0|download1_s1_translator|read_latency_shift_reg~0_combout ),
	.cp_valid(\mm_interconnect_0|cpu_data_master_agent|cp_valid~0_combout ),
	.W_debug_mode(\cpu|cpu|W_debug_mode~q ),
	.read_latency_shift_reg_0(\mm_interconnect_0|camstate1_s1_translator|read_latency_shift_reg[0]~q ),
	.WideOr1(\mm_interconnect_0|rsp_mux|WideOr1~0_combout ),
	.WideOr11(\mm_interconnect_0|rsp_mux|WideOr1~1_combout ),
	.src0_valid(\mm_interconnect_0|rsp_demux_002|src0_valid~0_combout ),
	.src0_valid1(\mm_interconnect_0|rsp_demux_003|src0_valid~0_combout ),
	.read_latency_shift_reg_01(\mm_interconnect_0|jtag_uart_avalon_jtag_slave_translator|read_latency_shift_reg[0]~q ),
	.WideOr12(\mm_interconnect_0|rsp_mux|WideOr1~3_combout ),
	.WideOr13(\mm_interconnect_0|rsp_mux|WideOr1~combout ),
	.Equal21(\mm_interconnect_0|router|Equal2~2_combout ),
	.wait_latency_counter_06(\mm_interconnect_0|sys_clk_timer_s1_translator|wait_latency_counter[0]~q ),
	.mem_used_14(\mm_interconnect_0|sys_clk_timer_s1_agent_rsp_fifo|mem_used[1]~q ),
	.wait_latency_counter_15(\mm_interconnect_0|sys_clk_timer_s1_translator|wait_latency_counter[1]~q ),
	.mem_used_15(\mm_interconnect_0|onchip_mem_s1_agent_rsp_fifo|mem_used[1]~q ),
	.saved_grant_0(\mm_interconnect_0|cmd_mux_003|saved_grant[0]~q ),
	.always11(\mm_interconnect_0|router|always1~2_combout ),
	.av_waitrequest(\jtag_uart|av_waitrequest~q ),
	.mem_used_16(\mm_interconnect_0|jtag_uart_avalon_jtag_slave_agent_rsp_fifo|mem_used[1]~q ),
	.av_waitrequest1(\jtag_uart|av_waitrequest~0_combout ),
	.saved_grant_01(\mm_interconnect_0|cmd_mux_002|saved_grant[0]~q ),
	.waitrequest(\cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|the_first_nios2_system_cpu_cpu_nios2_ocimem|waitrequest~q ),
	.mem_used_17(\mm_interconnect_0|cpu_debug_mem_slave_agent_rsp_fifo|mem_used[1]~q ),
	.cpu_data_master_waitrequest(\mm_interconnect_0|cpu_data_master_translator|av_waitrequest~0_combout ),
	.i_read(\cpu|cpu|i_read~q ),
	.ic_fill_tag_5(\cpu|cpu|ic_fill_tag[5]~q ),
	.ic_fill_tag_4(\cpu|cpu|ic_fill_tag[4]~q ),
	.ic_fill_tag_3(\cpu|cpu|ic_fill_tag[3]~q ),
	.ic_fill_tag_2(\cpu|cpu|ic_fill_tag[2]~q ),
	.ic_fill_tag_1(\cpu|cpu|ic_fill_tag[1]~q ),
	.ic_fill_tag_0(\cpu|cpu|ic_fill_tag[0]~q ),
	.WideOr14(\mm_interconnect_0|cmd_mux_002|WideOr1~combout ),
	.mem(\mm_interconnect_0|cpu_debug_mem_slave_agent_rsp_fifo|mem~0_combout ),
	.WideOr15(\mm_interconnect_0|cmd_mux_003|WideOr1~combout ),
	.ien_AE(\jtag_uart|ien_AE~q ),
	.av_readdata_9(\jtag_uart|av_readdata[9]~combout ),
	.ien_AF(\jtag_uart|ien_AF~q ),
	.av_readdata_8(\jtag_uart|av_readdata[8]~0_combout ),
	.src_payload(\mm_interconnect_0|cmd_mux_002|src_payload~0_combout ),
	.ic_fill_ap_offset_0(\cpu|cpu|ic_fill_ap_offset[0]~q ),
	.src_data_38(\mm_interconnect_0|cmd_mux_002|src_data[38]~combout ),
	.ic_fill_line_0(\cpu|cpu|ic_fill_line[0]~q ),
	.src_data_41(\mm_interconnect_0|cmd_mux_002|src_data[41]~combout ),
	.ic_fill_ap_offset_2(\cpu|cpu|ic_fill_ap_offset[2]~q ),
	.src_data_40(\mm_interconnect_0|cmd_mux_002|src_data[40]~combout ),
	.ic_fill_ap_offset_1(\cpu|cpu|ic_fill_ap_offset[1]~q ),
	.src_data_39(\mm_interconnect_0|cmd_mux_002|src_data[39]~combout ),
	.ic_fill_line_5(\cpu|cpu|ic_fill_line[5]~q ),
	.src_data_46(\mm_interconnect_0|cmd_mux_002|src_data[46]~combout ),
	.ic_fill_line_4(\cpu|cpu|ic_fill_line[4]~q ),
	.src_data_45(\mm_interconnect_0|cmd_mux_002|src_data[45]~combout ),
	.ic_fill_line_3(\cpu|cpu|ic_fill_line[3]~q ),
	.src_data_44(\mm_interconnect_0|cmd_mux_002|src_data[44]~combout ),
	.ic_fill_line_2(\cpu|cpu|ic_fill_line[2]~q ),
	.src_data_43(\mm_interconnect_0|cmd_mux_002|src_data[43]~combout ),
	.ic_fill_line_1(\cpu|cpu|ic_fill_line[1]~q ),
	.src_data_42(\mm_interconnect_0|cmd_mux_002|src_data[42]~combout ),
	.src_payload1(\mm_interconnect_0|cmd_mux_002|src_payload~1_combout ),
	.save_dest_id(\mm_interconnect_0|cpu_instruction_master_limiter|save_dest_id~0_combout ),
	.WideOr0(\mm_interconnect_0|cmd_demux_001|WideOr0~0_combout ),
	.nonposted_cmd_accepted(\mm_interconnect_0|cpu_instruction_master_limiter|nonposted_cmd_accepted~combout ),
	.suppress_change_dest_id(\mm_interconnect_0|cpu_instruction_master_limiter|suppress_change_dest_id~0_combout ),
	.b_full(\jtag_uart|the_first_nios2_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|b_full~q ),
	.src_data_0(\mm_interconnect_0|rsp_mux|src_data[0]~combout ),
	.b_full1(\jtag_uart|the_first_nios2_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|b_full~q ),
	.b_non_empty(\jtag_uart|the_first_nios2_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|b_non_empty~q ),
	.read_0(\jtag_uart|read_0~q ),
	.counter_reg_bit_0(\jtag_uart|the_first_nios2_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[0]~q ),
	.src_payload2(\mm_interconnect_0|rsp_mux|src_payload~0_combout ),
	.src_data_1(\mm_interconnect_0|rsp_mux|src_data[1]~combout ),
	.src_data_2(\mm_interconnect_0|rsp_mux|src_data[2]~combout ),
	.src_data_3(\mm_interconnect_0|rsp_mux|src_data[3]~combout ),
	.src_payload3(\mm_interconnect_0|rsp_mux|src_payload~3_combout ),
	.src_payload4(\mm_interconnect_0|rsp_mux|src_payload~7_combout ),
	.src_payload5(\mm_interconnect_0|rsp_mux|src_payload~12_combout ),
	.src_payload6(\mm_interconnect_0|rsp_mux|src_payload~15_combout ),
	.src_payload7(\mm_interconnect_0|cmd_mux_002|src_payload~2_combout ),
	.A_mem_byte_en_0(\cpu|cpu|A_mem_byte_en[0]~q ),
	.src_data_32(\mm_interconnect_0|cmd_mux_002|src_data[32]~combout ),
	.counter_reg_bit_1(\jtag_uart|the_first_nios2_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[1]~q ),
	.counter_reg_bit_4(\jtag_uart|the_first_nios2_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[4]~q ),
	.counter_reg_bit_3(\jtag_uart|the_first_nios2_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[3]~q ),
	.counter_reg_bit_2(\jtag_uart|the_first_nios2_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[2]~q ),
	.counter_reg_bit_5(\jtag_uart|the_first_nios2_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[5]~q ),
	.av_readdata_pre_221(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[22]~q ),
	.src_payload8(\mm_interconnect_0|rsp_mux|src_payload~16_combout ),
	.av_readdata_pre_23(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[23]~q ),
	.src_payload9(\mm_interconnect_0|rsp_mux|src_payload~17_combout ),
	.av_readdata_pre_24(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[24]~q ),
	.src_payload10(\mm_interconnect_0|rsp_mux|src_payload~18_combout ),
	.av_readdata_pre_25(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[25]~q ),
	.src_payload11(\mm_interconnect_0|rsp_mux|src_payload~19_combout ),
	.av_readdata_pre_31(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[31]~q ),
	.src_payload12(\mm_interconnect_0|rsp_mux|src_payload~20_combout ),
	.av_readdata_pre_21(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[21]~q ),
	.src_payload13(\mm_interconnect_0|rsp_mux|src_payload~21_combout ),
	.src_payload14(\mm_interconnect_0|rsp_mux|src_payload~22_combout ),
	.av_readdata_pre_11(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[11]~q ),
	.src_payload15(\mm_interconnect_0|rsp_mux|src_payload~23_combout ),
	.src_payload16(\mm_interconnect_0|rsp_mux|src_payload~24_combout ),
	.av_readdata_pre_28(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[28]~q ),
	.src_payload17(\mm_interconnect_0|rsp_mux|src_payload~25_combout ),
	.av_readdata_pre_10(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[10]~q ),
	.src_payload18(\mm_interconnect_0|rsp_mux|src_payload~26_combout ),
	.src_payload19(\mm_interconnect_0|rsp_mux|src_payload~27_combout ),
	.av_readdata_pre_27(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[27]~q ),
	.src_payload20(\mm_interconnect_0|rsp_mux|src_payload~28_combout ),
	.av_readdata_pre_8(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[8]~q ),
	.src_payload21(\mm_interconnect_0|rsp_mux|src_payload~29_combout ),
	.src_payload22(\mm_interconnect_0|rsp_mux|src_payload~30_combout ),
	.av_readdata_pre_9(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[9]~q ),
	.src_payload23(\mm_interconnect_0|rsp_mux|src_payload~31_combout ),
	.src_payload24(\mm_interconnect_0|rsp_mux|src_payload~32_combout ),
	.av_readdata_pre_26(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[26]~q ),
	.src_payload25(\mm_interconnect_0|rsp_mux|src_payload~33_combout ),
	.av_readdata_pre_201(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[20]~q ),
	.src_payload26(\mm_interconnect_0|rsp_mux|src_payload~34_combout ),
	.av_readdata_pre_191(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[19]~q ),
	.src_payload27(\mm_interconnect_0|rsp_mux|src_payload~35_combout ),
	.av_readdata_pre_17(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[17]~q ),
	.src_payload28(\mm_interconnect_0|rsp_mux|src_payload~36_combout ),
	.src_payload29(\mm_interconnect_0|rsp_mux|src_payload~37_combout ),
	.av_readdata_pre_30(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[30]~q ),
	.src_payload30(\mm_interconnect_0|rsp_mux|src_payload~38_combout ),
	.av_readdata_pre_18(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[18]~q ),
	.src_payload31(\mm_interconnect_0|rsp_mux|src_payload~39_combout ),
	.src_payload32(\mm_interconnect_0|rsp_mux|src_payload~40_combout ),
	.av_readdata_pre_16(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[16]~q ),
	.src_payload33(\mm_interconnect_0|rsp_mux|src_payload~41_combout ),
	.src_payload34(\mm_interconnect_0|rsp_mux|src_payload~42_combout ),
	.av_readdata_pre_15(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[15]~q ),
	.src_payload35(\mm_interconnect_0|rsp_mux|src_payload~43_combout ),
	.src_payload36(\mm_interconnect_0|rsp_mux|src_payload~44_combout ),
	.av_readdata_pre_12(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[12]~q ),
	.src_payload37(\mm_interconnect_0|rsp_mux|src_payload~45_combout ),
	.src_payload38(\mm_interconnect_0|rsp_mux|src_payload~46_combout ),
	.av_readdata_pre_13(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[13]~q ),
	.src_payload39(\mm_interconnect_0|rsp_mux|src_payload~47_combout ),
	.src_payload40(\mm_interconnect_0|rsp_mux|src_payload~48_combout ),
	.av_readdata_pre_14(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[14]~q ),
	.src_payload41(\mm_interconnect_0|rsp_mux|src_payload~49_combout ),
	.src_payload42(\mm_interconnect_0|rsp_mux|src_payload~50_combout ),
	.av_readdata_pre_29(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[29]~q ),
	.src_payload43(\mm_interconnect_0|rsp_mux|src_payload~51_combout ),
	.src_payload44(\mm_interconnect_0|cmd_mux_003|src_payload~0_combout ),
	.src_data_381(\mm_interconnect_0|cmd_mux_003|src_data[38]~combout ),
	.src_data_391(\mm_interconnect_0|cmd_mux_003|src_data[39]~combout ),
	.src_data_401(\mm_interconnect_0|cmd_mux_003|src_data[40]~combout ),
	.src_data_411(\mm_interconnect_0|cmd_mux_003|src_data[41]~combout ),
	.src_data_421(\mm_interconnect_0|cmd_mux_003|src_data[42]~combout ),
	.src_data_431(\mm_interconnect_0|cmd_mux_003|src_data[43]~combout ),
	.src_data_441(\mm_interconnect_0|cmd_mux_003|src_data[44]~combout ),
	.src_data_451(\mm_interconnect_0|cmd_mux_003|src_data[45]~combout ),
	.src_data_461(\mm_interconnect_0|cmd_mux_003|src_data[46]~combout ),
	.src_data_47(\mm_interconnect_0|cmd_mux_003|src_data[47]~combout ),
	.src_data_48(\mm_interconnect_0|cmd_mux_003|src_data[48]~combout ),
	.src_data_49(\mm_interconnect_0|cmd_mux_003|src_data[49]~combout ),
	.src_data_50(\mm_interconnect_0|cmd_mux_003|src_data[50]~combout ),
	.src_data_321(\mm_interconnect_0|cmd_mux_003|src_data[32]~combout ),
	.readdata_09(\sys_clk_timer|readdata[0]~q ),
	.src_payload45(\mm_interconnect_0|cmd_mux_002|src_payload~3_combout ),
	.A_st_data_16(\cpu|cpu|A_st_data[16]~q ),
	.src_payload46(\mm_interconnect_0|cmd_mux_002|src_payload~4_combout ),
	.WideOr16(\mm_interconnect_0|rsp_mux_001|WideOr1~combout ),
	.src_payload47(\mm_interconnect_0|cmd_mux_003|src_payload~1_combout ),
	.readdata_110(\sys_clk_timer|readdata[1]~q ),
	.src_payload48(\mm_interconnect_0|cmd_mux_003|src_payload~2_combout ),
	.readdata_210(\sys_clk_timer|readdata[2]~q ),
	.src_payload49(\mm_interconnect_0|cmd_mux_003|src_payload~3_combout ),
	.readdata_37(\sys_clk_timer|readdata[3]~q ),
	.readdata_45(\sys_clk_timer|readdata[4]~q ),
	.src_payload50(\mm_interconnect_0|cmd_mux_003|src_payload~4_combout ),
	.src_payload51(\mm_interconnect_0|cmd_mux_003|src_payload~5_combout ),
	.readdata_55(\sys_clk_timer|readdata[5]~q ),
	.src_payload52(\mm_interconnect_0|cmd_mux_003|src_payload~6_combout ),
	.readdata_63(\sys_clk_timer|readdata[6]~q ),
	.src_payload53(\mm_interconnect_0|cmd_mux_003|src_payload~7_combout ),
	.readdata_71(\sys_clk_timer|readdata[7]~q ),
	.A_st_data_22(\cpu|cpu|A_st_data[22]~q ),
	.src_payload54(\mm_interconnect_0|cmd_mux_003|src_payload~8_combout ),
	.A_mem_byte_en_2(\cpu|cpu|A_mem_byte_en[2]~q ),
	.src_data_34(\mm_interconnect_0|cmd_mux_003|src_data[34]~combout ),
	.A_st_data_23(\cpu|cpu|A_st_data[23]~q ),
	.src_payload55(\mm_interconnect_0|cmd_mux_003|src_payload~9_combout ),
	.A_st_data_24(\cpu|cpu|A_st_data[24]~q ),
	.src_payload56(\mm_interconnect_0|cmd_mux_003|src_payload~10_combout ),
	.A_mem_byte_en_3(\cpu|cpu|A_mem_byte_en[3]~q ),
	.src_data_35(\mm_interconnect_0|cmd_mux_003|src_data[35]~combout ),
	.A_st_data_25(\cpu|cpu|A_st_data[25]~q ),
	.src_payload57(\mm_interconnect_0|cmd_mux_003|src_payload~11_combout ),
	.A_st_data_31(\cpu|cpu|A_st_data[31]~q ),
	.src_payload58(\mm_interconnect_0|cmd_mux_003|src_payload~12_combout ),
	.A_st_data_21(\cpu|cpu|A_st_data[21]~q ),
	.src_payload59(\mm_interconnect_0|cmd_mux_003|src_payload~13_combout ),
	.A_st_data_11(\cpu|cpu|A_st_data[11]~q ),
	.src_payload60(\mm_interconnect_0|cmd_mux_003|src_payload~14_combout ),
	.A_mem_byte_en_1(\cpu|cpu|A_mem_byte_en[1]~q ),
	.src_data_33(\mm_interconnect_0|cmd_mux_003|src_data[33]~combout ),
	.readdata_112(\sys_clk_timer|readdata[11]~q ),
	.A_st_data_28(\cpu|cpu|A_st_data[28]~q ),
	.src_payload61(\mm_interconnect_0|cmd_mux_003|src_payload~15_combout ),
	.A_st_data_10(\cpu|cpu|A_st_data[10]~q ),
	.src_payload62(\mm_interconnect_0|cmd_mux_003|src_payload~16_combout ),
	.ac(\jtag_uart|ac~q ),
	.readdata_101(\sys_clk_timer|readdata[10]~q ),
	.A_st_data_27(\cpu|cpu|A_st_data[27]~q ),
	.src_payload63(\mm_interconnect_0|cmd_mux_003|src_payload~17_combout ),
	.A_st_data_8(\cpu|cpu|A_st_data[8]~q ),
	.src_payload64(\mm_interconnect_0|cmd_mux_003|src_payload~18_combout ),
	.readdata_81(\sys_clk_timer|readdata[8]~q ),
	.A_st_data_9(\cpu|cpu|A_st_data[9]~q ),
	.src_payload65(\mm_interconnect_0|cmd_mux_003|src_payload~19_combout ),
	.readdata_91(\sys_clk_timer|readdata[9]~q ),
	.A_st_data_26(\cpu|cpu|A_st_data[26]~q ),
	.src_payload66(\mm_interconnect_0|cmd_mux_003|src_payload~20_combout ),
	.A_st_data_20(\cpu|cpu|A_st_data[20]~q ),
	.src_payload67(\mm_interconnect_0|cmd_mux_003|src_payload~21_combout ),
	.A_st_data_19(\cpu|cpu|A_st_data[19]~q ),
	.src_payload68(\mm_interconnect_0|cmd_mux_003|src_payload~22_combout ),
	.A_st_data_17(\cpu|cpu|A_st_data[17]~q ),
	.src_payload69(\mm_interconnect_0|cmd_mux_003|src_payload~23_combout ),
	.A_st_data_30(\cpu|cpu|A_st_data[30]~q ),
	.src_payload70(\mm_interconnect_0|cmd_mux_003|src_payload~24_combout ),
	.A_st_data_18(\cpu|cpu|A_st_data[18]~q ),
	.src_payload71(\mm_interconnect_0|cmd_mux_003|src_payload~25_combout ),
	.src_payload72(\mm_interconnect_0|cmd_mux_003|src_payload~26_combout ),
	.A_st_data_15(\cpu|cpu|A_st_data[15]~q ),
	.src_payload73(\mm_interconnect_0|cmd_mux_003|src_payload~27_combout ),
	.rvalid(\jtag_uart|rvalid~q ),
	.readdata_152(\sys_clk_timer|readdata[15]~q ),
	.A_st_data_12(\cpu|cpu|A_st_data[12]~q ),
	.src_payload74(\mm_interconnect_0|cmd_mux_003|src_payload~28_combout ),
	.readdata_122(\sys_clk_timer|readdata[12]~q ),
	.A_st_data_13(\cpu|cpu|A_st_data[13]~q ),
	.src_payload75(\mm_interconnect_0|cmd_mux_003|src_payload~29_combout ),
	.readdata_132(\sys_clk_timer|readdata[13]~q ),
	.A_st_data_14(\cpu|cpu|A_st_data[14]~q ),
	.src_payload76(\mm_interconnect_0|cmd_mux_003|src_payload~30_combout ),
	.woverflow(\jtag_uart|woverflow~q ),
	.readdata_142(\sys_clk_timer|readdata[14]~q ),
	.A_st_data_29(\cpu|cpu|A_st_data[29]~q ),
	.src_payload77(\mm_interconnect_0|cmd_mux_003|src_payload~31_combout ),
	.src_data_26(\mm_interconnect_0|rsp_mux_001|src_data[26]~combout ),
	.src_data_25(\mm_interconnect_0|rsp_mux_001|src_data[25]~combout ),
	.src_data_24(\mm_interconnect_0|rsp_mux_001|src_data[24]~combout ),
	.src_data_23(\mm_interconnect_0|rsp_mux_001|src_data[23]~combout ),
	.src_data_22(\mm_interconnect_0|rsp_mux_001|src_data[22]~combout ),
	.src_data_11(\mm_interconnect_0|rsp_mux_001|src_data[1]~combout ),
	.src_data_01(\mm_interconnect_0|rsp_mux_001|src_data[0]~combout ),
	.src_data_21(\mm_interconnect_0|rsp_mux_001|src_data[2]~combout ),
	.src_data_31(\mm_interconnect_0|rsp_mux_001|src_data[3]~combout ),
	.src_data_4(\mm_interconnect_0|rsp_mux_001|src_data[4]~combout ),
	.src_data_5(\mm_interconnect_0|rsp_mux_001|src_data[5]~combout ),
	.src_data_28(\mm_interconnect_0|rsp_mux_001|src_data[28]~combout ),
	.src_data_311(\mm_interconnect_0|rsp_mux_001|src_data[31]~combout ),
	.src_data_27(\mm_interconnect_0|rsp_mux_001|src_data[27]~combout ),
	.src_data_29(\mm_interconnect_0|rsp_mux_001|src_data[29]~combout ),
	.src_data_30(\mm_interconnect_0|rsp_mux_001|src_data[30]~combout ),
	.src_data_111(\mm_interconnect_0|rsp_mux_001|src_data[11]~combout ),
	.src_data_12(\mm_interconnect_0|rsp_mux_001|src_data[12]~combout ),
	.src_data_13(\mm_interconnect_0|rsp_mux_001|src_data[13]~combout ),
	.src_data_14(\mm_interconnect_0|rsp_mux_001|src_data[14]~combout ),
	.src_data_15(\mm_interconnect_0|rsp_mux_001|src_data[15]~combout ),
	.src_data_16(\mm_interconnect_0|rsp_mux_001|src_data[16]~combout ),
	.src_payload78(\mm_interconnect_0|cmd_mux_002|src_payload~5_combout ),
	.src_data_9(\mm_interconnect_0|rsp_mux_001|src_data[9]~combout ),
	.src_data_211(\mm_interconnect_0|rsp_mux_001|src_data[21]~combout ),
	.src_data_6(\mm_interconnect_0|rsp_mux_001|src_data[6]~combout ),
	.src_data_8(\mm_interconnect_0|rsp_mux_001|src_data[8]~combout ),
	.src_data_17(\mm_interconnect_0|rsp_mux_001|src_data[17]~combout ),
	.src_data_18(\mm_interconnect_0|rsp_mux_001|src_data[18]~combout ),
	.src_data_10(\mm_interconnect_0|rsp_mux_001|src_data[10]~combout ),
	.src_data_7(\mm_interconnect_0|rsp_mux_001|src_data[7]~combout ),
	.src_data_20(\mm_interconnect_0|rsp_mux_001|src_data[20]~combout ),
	.src_data_19(\mm_interconnect_0|rsp_mux_001|src_data[19]~combout ),
	.src_payload79(\mm_interconnect_0|cmd_mux_002|src_payload~6_combout ),
	.src_data_341(\mm_interconnect_0|cmd_mux_002|src_data[34]~combout ),
	.src_payload80(\mm_interconnect_0|cmd_mux_002|src_payload~7_combout ),
	.src_payload81(\mm_interconnect_0|cmd_mux_002|src_payload~8_combout ),
	.src_payload82(\mm_interconnect_0|cmd_mux_002|src_payload~9_combout ),
	.src_payload83(\mm_interconnect_0|cmd_mux_002|src_payload~10_combout ),
	.src_payload84(\mm_interconnect_0|cmd_mux_002|src_payload~11_combout ),
	.src_payload85(\mm_interconnect_0|cmd_mux_002|src_payload~12_combout ),
	.src_payload86(\mm_interconnect_0|cmd_mux_002|src_payload~13_combout ),
	.src_payload87(\mm_interconnect_0|cmd_mux_002|src_payload~14_combout ),
	.src_payload88(\mm_interconnect_0|cmd_mux_002|src_payload~15_combout ),
	.src_data_351(\mm_interconnect_0|cmd_mux_002|src_data[35]~combout ),
	.src_payload89(\mm_interconnect_0|cmd_mux_002|src_payload~16_combout ),
	.src_payload90(\mm_interconnect_0|cmd_mux_002|src_payload~17_combout ),
	.src_payload91(\mm_interconnect_0|cmd_mux_002|src_payload~18_combout ),
	.src_payload92(\mm_interconnect_0|cmd_mux_002|src_payload~19_combout ),
	.src_payload93(\mm_interconnect_0|cmd_mux_002|src_payload~20_combout ),
	.src_payload94(\mm_interconnect_0|cmd_mux_002|src_payload~21_combout ),
	.src_payload95(\mm_interconnect_0|cmd_mux_002|src_payload~22_combout ),
	.src_data_331(\mm_interconnect_0|cmd_mux_002|src_data[33]~combout ),
	.src_payload96(\mm_interconnect_0|cmd_mux_002|src_payload~23_combout ),
	.src_payload97(\mm_interconnect_0|cmd_mux_002|src_payload~24_combout ),
	.src_payload98(\mm_interconnect_0|cmd_mux_002|src_payload~25_combout ),
	.src_payload99(\mm_interconnect_0|cmd_mux_002|src_payload~26_combout ),
	.src_payload100(\mm_interconnect_0|cmd_mux_002|src_payload~27_combout ),
	.src_payload101(\mm_interconnect_0|cmd_mux_002|src_payload~28_combout ),
	.src_payload102(\mm_interconnect_0|cmd_mux_002|src_payload~29_combout ),
	.src_payload103(\mm_interconnect_0|cmd_mux_002|src_payload~30_combout ),
	.src_payload104(\mm_interconnect_0|cmd_mux_002|src_payload~31_combout ),
	.src_payload105(\mm_interconnect_0|cmd_mux_002|src_payload~32_combout ),
	.GND_port(\~GND~combout ),
	.clk_clk(\clk_clk~input_o ));

first_nios2_system_first_nios2_system_tenOut1_1 tenout2(
	.readdata_0(\tenout2|readdata[0]~q ),
	.readdata_1(\tenout2|readdata[1]~q ),
	.readdata_2(\tenout2|readdata[2]~q ),
	.readdata_3(\tenout2|readdata[3]~q ),
	.Equal0(\camdata1|Equal0~0_combout ),
	.r_sync_rst(\rst_controller|r_sync_rst~q ),
	.clk_clk(\clk_clk~input_o ),
	.tenout2_external_connection_export_0(\tenout2_external_connection_export[0]~input_o ),
	.tenout2_external_connection_export_1(\tenout2_external_connection_export[1]~input_o ),
	.tenout2_external_connection_export_2(\tenout2_external_connection_export[2]~input_o ),
	.tenout2_external_connection_export_3(\tenout2_external_connection_export[3]~input_o ));

first_nios2_system_first_nios2_system_tenOut1 tenout1(
	.readdata_0(\tenout1|readdata[0]~q ),
	.readdata_1(\tenout1|readdata[1]~q ),
	.readdata_2(\tenout1|readdata[2]~q ),
	.readdata_3(\tenout1|readdata[3]~q ),
	.Equal0(\camdata1|Equal0~0_combout ),
	.r_sync_rst(\rst_controller|r_sync_rst~q ),
	.clk_clk(\clk_clk~input_o ),
	.tenout1_external_connection_export_0(\tenout1_external_connection_export[0]~input_o ),
	.tenout1_external_connection_export_1(\tenout1_external_connection_export[1]~input_o ),
	.tenout1_external_connection_export_2(\tenout1_external_connection_export[2]~input_o ),
	.tenout1_external_connection_export_3(\tenout1_external_connection_export[3]~input_o ));

first_nios2_system_altera_reset_controller rst_controller(
	.r_sync_rst1(\rst_controller|r_sync_rst~q ),
	.r_early_rst1(\rst_controller|r_early_rst~q ),
	.altera_reset_synchronizer_int_chain_1(\rst_controller|alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain[1]~0_combout ),
	.clk_clk(\clk_clk~input_o ),
	.reset_reset_n(\reset_reset_n~input_o ));

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_1[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_1[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_1[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_1[3] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~3_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~5_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~6_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~5_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0 .lut_mask = 64'hFEFEFEFEFEFEFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\altera_internal_jtag~TDIUTAP ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1 .lut_mask = 64'hEDDEFFFFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2 .lut_mask = 64'h7FBFFFFFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\altera_internal_jtag~TDIUTAP ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3 .lut_mask = 64'hFFFFB77BFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~5_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~6_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~3 .lut_mask = 64'h4747474747474747;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~3 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~14 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~14 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~14 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~14 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~4 .lut_mask = 64'hFFFFEFFFFFFFFFEF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~4 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~5 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~14_combout ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~4_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~5 .lut_mask = 64'hFFF7FFFFFFF7FFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~5 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~7_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~6_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~6 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~6 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~6 .lut_mask = 64'h4747474747474747;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~6 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~5 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~5 .lut_mask = 64'h2727272727272727;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~5 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~6 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~14_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~6 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~6 .lut_mask = 64'hFFFFFFFF7FFFF7FF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~6 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~7 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~7 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~7 .lut_mask = 64'h2727272727272727;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~7 .shared_arith = "off";

assign \clk_clk~input_o  = clk_clk;

assign \camstate2_external_connection_export[0]~input_o  = camstate2_external_connection_export[0];

assign \tenout1_external_connection_export[0]~input_o  = tenout1_external_connection_export[0];

assign \tenout2_external_connection_export[0]~input_o  = tenout2_external_connection_export[0];

assign \camstate1_external_connection_export[0]~input_o  = camstate1_external_connection_export[0];

assign \rtd2_external_connection_export~input_o  = rtd2_external_connection_export;

assign \rtd1_external_connection_export~input_o  = rtd1_external_connection_export;

assign \camdata1_external_connection_export[0]~input_o  = camdata1_external_connection_export[0];

assign \camdata2_external_connection_export[0]~input_o  = camdata2_external_connection_export[0];

assign \reset_reset_n~input_o  = reset_reset_n;

assign \tenout2_external_connection_export[1]~input_o  = tenout2_external_connection_export[1];

assign \camdata1_external_connection_export[1]~input_o  = camdata1_external_connection_export[1];

assign \camstate2_external_connection_export[1]~input_o  = camstate2_external_connection_export[1];

assign \camdata2_external_connection_export[1]~input_o  = camdata2_external_connection_export[1];

assign \camstate1_external_connection_export[1]~input_o  = camstate1_external_connection_export[1];

assign \tenout1_external_connection_export[1]~input_o  = tenout1_external_connection_export[1];

assign \tenout2_external_connection_export[2]~input_o  = tenout2_external_connection_export[2];

assign \camdata1_external_connection_export[2]~input_o  = camdata1_external_connection_export[2];

assign \camstate2_external_connection_export[2]~input_o  = camstate2_external_connection_export[2];

assign \camdata2_external_connection_export[2]~input_o  = camdata2_external_connection_export[2];

assign \camstate1_external_connection_export[2]~input_o  = camstate1_external_connection_export[2];

assign \tenout1_external_connection_export[2]~input_o  = tenout1_external_connection_export[2];

assign \camdata2_external_connection_export[3]~input_o  = camdata2_external_connection_export[3];

assign \tenout2_external_connection_export[3]~input_o  = tenout2_external_connection_export[3];

assign \camdata1_external_connection_export[3]~input_o  = camdata1_external_connection_export[3];

assign \tenout1_external_connection_export[3]~input_o  = tenout1_external_connection_export[3];

assign \camstate1_external_connection_export[3]~input_o  = camstate1_external_connection_export[3];

assign \camstate2_external_connection_export[3]~input_o  = camstate2_external_connection_export[3];

assign \camdata1_external_connection_export[4]~input_o  = camdata1_external_connection_export[4];

assign \camdata2_external_connection_export[4]~input_o  = camdata2_external_connection_export[4];

assign \camstate1_external_connection_export[4]~input_o  = camstate1_external_connection_export[4];

assign \camstate2_external_connection_export[4]~input_o  = camstate2_external_connection_export[4];

assign \camdata1_external_connection_export[5]~input_o  = camdata1_external_connection_export[5];

assign \camdata2_external_connection_export[5]~input_o  = camdata2_external_connection_export[5];

assign \camstate1_external_connection_export[5]~input_o  = camstate1_external_connection_export[5];

assign \camstate2_external_connection_export[5]~input_o  = camstate2_external_connection_export[5];

assign \camdata1_external_connection_export[6]~input_o  = camdata1_external_connection_export[6];

assign \camdata2_external_connection_export[6]~input_o  = camdata2_external_connection_export[6];

assign download1_external_connection_export = \download1|data_out~q ;

assign download2_external_connection_export = \download2|data_out~q ;

assign hex1_external_connection_export[0] = \hex1|data_out[0]~q ;

assign hex1_external_connection_export[1] = \hex1|data_out[1]~q ;

assign hex1_external_connection_export[2] = \hex1|data_out[2]~q ;

assign hex1_external_connection_export[3] = \hex1|data_out[3]~q ;

assign hex1_external_connection_export[4] = \hex1|data_out[4]~q ;

assign hex1_external_connection_export[5] = \hex1|data_out[5]~q ;

assign hex1_external_connection_export[6] = \hex1|data_out[6]~q ;

assign hex2_external_connection_export[0] = \hex2|data_out[0]~q ;

assign hex2_external_connection_export[1] = \hex2|data_out[1]~q ;

assign hex2_external_connection_export[2] = \hex2|data_out[2]~q ;

assign hex2_external_connection_export[3] = \hex2|data_out[3]~q ;

assign hex2_external_connection_export[4] = \hex2|data_out[4]~q ;

assign hex2_external_connection_export[5] = \hex2|data_out[5]~q ;

assign hex2_external_connection_export[6] = \hex2|data_out[6]~q ;

assign leds_external_connection_export[0] = \leds|data_out[0]~q ;

assign leds_external_connection_export[1] = \leds|data_out[1]~q ;

assign leds_external_connection_export[2] = \leds|data_out[2]~q ;

assign leds_external_connection_export[3] = \leds|data_out[3]~q ;

assign leds_external_connection_export[4] = \leds|data_out[4]~q ;

assign leds_external_connection_export[5] = \leds|data_out[5]~q ;

assign leds_external_connection_export[6] = \leds|data_out[6]~q ;

assign leds_external_connection_export[7] = \leds|data_out[7]~q ;

assign start_external_connection_export = \start|data_out~q ;

assign altera_reserved_tdo = \altera_internal_jtag~TDO ;

assign \altera_reserved_tms~input_o  = altera_reserved_tms;

assign \altera_reserved_tck~input_o  = altera_reserved_tck;

assign \altera_reserved_tdi~input_o  = altera_reserved_tdi;

cyclonev_jtag altera_internal_jtag(
	.tms(\altera_reserved_tms~input_o ),
	.tck(\altera_reserved_tck~input_o ),
	.tdi(\altera_reserved_tdi~input_o ),
	.tdoutap(gnd),
	.tdouser(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~q ),
	.tdo(\altera_internal_jtag~TDO ),
	.tmsutap(\altera_internal_jtag~TMSUTAP ),
	.tckutap(\altera_internal_jtag~TCKUTAP ),
	.tdiutap(\altera_internal_jtag~TDIUTAP ),
	.shiftuser(),
	.clkdruser(),
	.updateuser(),
	.runidleuser(),
	.usr1user());

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2 .lut_mask = 64'h6666666666666666;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0 .lut_mask = 64'h9696969696969696;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0 .lut_mask = 64'hFFFBFFFBFFFBFFFB;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\altera_internal_jtag~TDIUTAP ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0 .lut_mask = 64'hFFFFFFEFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg .power_up = "low";

cyclonev_lcell_comb \~GND (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\~GND~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \~GND .extended_lut = "off";
defparam \~GND .lut_mask = 64'h0000000000000000;
defparam \~GND .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~8 (
	.dataa(!\rst_controller|alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain[1]~0_combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datac(!\~GND~combout ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.dataf(!\altera_internal_jtag~TDIUTAP ),
	.datag(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~8 .extended_lut = "on";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~8 .lut_mask = 64'hEFFEFAFCEFFEFAFC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~8 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~5 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~5 .lut_mask = 64'h96FFFFFF96FFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~5 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~5_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~6 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~6 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~6 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~6 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datad(!\cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_tck|ir_out[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4 .lut_mask = 64'h47FF47FF47FF47FF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4_combout ),
	.asdata(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg~3 .lut_mask = 64'hFFFFFFDFFFFFFFDF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg~3 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg~3_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~1 .lut_mask = 64'hFFFFFFACFFFFFFAC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~1 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2 .lut_mask = 64'hDF1FDF1FDF1FDF1F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~6_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~7 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~7 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~7 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~7 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~7_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~3 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~3 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~3_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0_combout ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0 .lut_mask = 64'hFDDFFFFFDFFDFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~1 .lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~1 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2 .lut_mask = 64'hCF5FFFFFCF5FFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~8_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~1 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~1 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~2 .lut_mask = 64'hEFFFEFFFEFFFEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~2 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~3 .lut_mask = 64'h2727272727272727;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~3 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8_combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~1_combout ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~2_combout ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~4 .lut_mask = 64'h6F9F9F6FFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~4 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~4_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0 .lut_mask = 64'hEFDFDFEFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~0 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~0 .lut_mask = 64'hF7FFFFFFF7FFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~1 .lut_mask = 64'hF7FFFFF7FFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~1 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0_combout ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~0_combout ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~2 .lut_mask = 64'h7FFFF7FFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~2_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datab(!\cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_tck|ir_out[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~0 .lut_mask = 64'hB77BFFFFB77BFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~0_combout ),
	.asdata(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[1] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datac(!\jtag_uart|first_nios2_system_jtag_uart_alt_jtag_atlantic|tdo~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0 .lut_mask = 64'hFF3F7F7FFF3F7F7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~5 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~5 .lut_mask = 64'hFFAAAAFFAAFFFFAA;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~5 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1 .lut_mask = 64'hFFFFFFDFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~1 .lut_mask = 64'hF7FFFFFFF7FFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~2 .lut_mask = 64'hEBBEBEEBBEEBEBBE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~0 .lut_mask = 64'hFBFEFEFBFEFBFBFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~4 .lut_mask = 64'hFFFFFEFFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~4 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~3 .lut_mask = 64'hAAFFFFAAAAFFFFAA;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~3 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5 .lut_mask = 64'hFFFFFEFFFFFFFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datac(!\altera_internal_jtag~TDIUTAP ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datag(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8 .extended_lut = "on";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8 .lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~2 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6 .lut_mask = 64'hDF8FDF8FDF8FDF8F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5_combout ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7 .lut_mask = 64'hD8FFFFFFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~3 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~3 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4 .lut_mask = 64'hFFFFFFFFDF8FFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~0 .lut_mask = 64'h6996699669966996;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~1 .lut_mask = 64'hF7B3FFFFF7B3FFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0_combout ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1 .lut_mask = 64'hFFFEFFFFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datad(!\jtag_uart|first_nios2_system_jtag_uart_alt_jtag_atlantic|tdo~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[1]~q ),
	.dataf(!\cpu|cpu|the_first_nios2_system_cpu_cpu_nios2_oci|the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0 (
	.dataa(!\altera_internal_jtag~TDIUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0 .lut_mask = 64'h4747474747474747;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3 (
	.dataa(!\altera_internal_jtag~TDIUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~0 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~0 .lut_mask = 64'hAAAAAAAAFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~1 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datae(gnd),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~4 .lut_mask = 64'h55AA55AAFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~4 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~5 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~5 .lut_mask = 64'hAA5555AAFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~5 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datac(gnd),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~2 .lut_mask = 64'h66999966FFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~3 .lut_mask = 64'h96696996FFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~3 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~1 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~2 .lut_mask = 64'hFFFFFBFEFFFFFBFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~2 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7 .lut_mask = 64'h9669699696696996;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9 .lut_mask = 64'h9669699696696996;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0_combout ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0 .lut_mask = 64'hDFFFFFFFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\altera_internal_jtag~TDIUTAP ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0 .lut_mask = 64'hFBFFFFFFFBFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~10 (
	.dataa(!\altera_internal_jtag~TDIUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~0_combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~1_combout ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9_combout ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~10 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~10 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~10 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~4 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~4 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~4_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~0_combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~1_combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7_combout ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~4_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5 .lut_mask = 64'hFFFFF9F6FFFFF9F6;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~0_combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~1_combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6 .lut_mask = 64'h27FFFFFF27FFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~4_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~0_combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~1_combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~2_combout ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~3 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~3 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~4_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3 .lut_mask = 64'h4747474747474747;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5 .lut_mask = 64'hFFFFFFFFFFFFBFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3_combout ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4_combout ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6 .lut_mask = 64'hFFFFFFFFFFFBFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~7 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0_combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1_combout ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2_combout ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~7 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~7 .lut_mask = 64'hFFFF7FFFFFFF7FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~7 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo (
	.clk(!\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo .power_up = "low";

cyclonev_lcell_comb \auto_hub|~GND (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|~GND~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|~GND .extended_lut = "off";
defparam \auto_hub|~GND .lut_mask = 64'h0000000000000000;
defparam \auto_hub|~GND .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell .shared_arith = "off";

endmodule

module first_nios2_system_altera_reset_controller (
	r_sync_rst1,
	r_early_rst1,
	altera_reset_synchronizer_int_chain_1,
	clk_clk,
	reset_reset_n)/* synthesis synthesis_greybox=1 */;
output 	r_sync_rst1;
output 	r_early_rst1;
output 	altera_reset_synchronizer_int_chain_1;
input 	clk_clk;
input 	reset_reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain_out~q ;
wire \alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ;
wire \altera_reset_synchronizer_int_chain[0]~q ;
wire \altera_reset_synchronizer_int_chain[1]~q ;
wire \altera_reset_synchronizer_int_chain[2]~q ;
wire \altera_reset_synchronizer_int_chain[3]~q ;
wire \altera_reset_synchronizer_int_chain[4]~0_combout ;
wire \altera_reset_synchronizer_int_chain[4]~q ;
wire \r_sync_rst_chain[3]~q ;
wire \r_sync_rst_chain~1_combout ;
wire \r_sync_rst_chain[2]~q ;
wire \r_sync_rst_chain~0_combout ;
wire \r_sync_rst_chain[1]~q ;
wire \WideOr0~0_combout ;
wire \always2~0_combout ;


first_nios2_system_altera_reset_synchronizer alt_rst_req_sync_uq1(
	.altera_reset_synchronizer_int_chain_out1(\alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.altera_reset_synchronizer_int_chain_1(altera_reset_synchronizer_int_chain_1),
	.clk(clk_clk));

first_nios2_system_altera_reset_synchronizer_1 alt_rst_sync_uq1(
	.altera_reset_synchronizer_int_chain_out1(\alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.clk(clk_clk),
	.reset_reset_n(reset_reset_n));

dffeas r_sync_rst(
	.clk(clk_clk),
	.d(\WideOr0~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(r_sync_rst1),
	.prn(vcc));
defparam r_sync_rst.is_wysiwyg = "true";
defparam r_sync_rst.power_up = "low";

dffeas r_early_rst(
	.clk(clk_clk),
	.d(\always2~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(r_early_rst1),
	.prn(vcc));
defparam r_early_rst.is_wysiwyg = "true";
defparam r_early_rst.power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[0] (
	.clk(clk_clk),
	.d(\alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[0]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[0] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[0] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[1] (
	.clk(clk_clk),
	.d(\altera_reset_synchronizer_int_chain[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[1]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[1] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[1] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[2] (
	.clk(clk_clk),
	.d(\altera_reset_synchronizer_int_chain[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[2]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[2] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[2] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[3] (
	.clk(clk_clk),
	.d(\altera_reset_synchronizer_int_chain[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[3]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[3] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[3] .power_up = "low";

cyclonev_lcell_comb \altera_reset_synchronizer_int_chain[4]~0 (
	.dataa(!\altera_reset_synchronizer_int_chain[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\altera_reset_synchronizer_int_chain[4]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \altera_reset_synchronizer_int_chain[4]~0 .extended_lut = "off";
defparam \altera_reset_synchronizer_int_chain[4]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \altera_reset_synchronizer_int_chain[4]~0 .shared_arith = "off";

dffeas \altera_reset_synchronizer_int_chain[4] (
	.clk(clk_clk),
	.d(\altera_reset_synchronizer_int_chain[4]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[4]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[4] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[4] .power_up = "low";

dffeas \r_sync_rst_chain[3] (
	.clk(clk_clk),
	.d(\altera_reset_synchronizer_int_chain[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\r_sync_rst_chain[3]~q ),
	.prn(vcc));
defparam \r_sync_rst_chain[3] .is_wysiwyg = "true";
defparam \r_sync_rst_chain[3] .power_up = "low";

cyclonev_lcell_comb \r_sync_rst_chain~1 (
	.dataa(!\altera_reset_synchronizer_int_chain[2]~q ),
	.datab(!\r_sync_rst_chain[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\r_sync_rst_chain~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \r_sync_rst_chain~1 .extended_lut = "off";
defparam \r_sync_rst_chain~1 .lut_mask = 64'h7777777777777777;
defparam \r_sync_rst_chain~1 .shared_arith = "off";

dffeas \r_sync_rst_chain[2] (
	.clk(clk_clk),
	.d(\r_sync_rst_chain~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\r_sync_rst_chain[2]~q ),
	.prn(vcc));
defparam \r_sync_rst_chain[2] .is_wysiwyg = "true";
defparam \r_sync_rst_chain[2] .power_up = "low";

cyclonev_lcell_comb \r_sync_rst_chain~0 (
	.dataa(!\altera_reset_synchronizer_int_chain[2]~q ),
	.datab(!\r_sync_rst_chain[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\r_sync_rst_chain~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \r_sync_rst_chain~0 .extended_lut = "off";
defparam \r_sync_rst_chain~0 .lut_mask = 64'h7777777777777777;
defparam \r_sync_rst_chain~0 .shared_arith = "off";

dffeas \r_sync_rst_chain[1] (
	.clk(clk_clk),
	.d(\r_sync_rst_chain~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\r_sync_rst_chain[1]~q ),
	.prn(vcc));
defparam \r_sync_rst_chain[1] .is_wysiwyg = "true";
defparam \r_sync_rst_chain[1] .power_up = "low";

cyclonev_lcell_comb \WideOr0~0 (
	.dataa(!r_sync_rst1),
	.datab(!\altera_reset_synchronizer_int_chain[4]~q ),
	.datac(!\r_sync_rst_chain[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~0 .extended_lut = "off";
defparam \WideOr0~0 .lut_mask = 64'hF7F7F7F7F7F7F7F7;
defparam \WideOr0~0 .shared_arith = "off";

cyclonev_lcell_comb \always2~0 (
	.dataa(!\r_sync_rst_chain[2]~q ),
	.datab(!\alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always2~0 .extended_lut = "off";
defparam \always2~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \always2~0 .shared_arith = "off";

endmodule

module first_nios2_system_altera_reset_synchronizer (
	altera_reset_synchronizer_int_chain_out1,
	altera_reset_synchronizer_int_chain_1,
	clk)/* synthesis synthesis_greybox=1 */;
output 	altera_reset_synchronizer_int_chain_out1;
output 	altera_reset_synchronizer_int_chain_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \altera_reset_synchronizer_int_chain[1]~q ;
wire \altera_reset_synchronizer_int_chain[0]~q ;


dffeas altera_reset_synchronizer_int_chain_out(
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(altera_reset_synchronizer_int_chain_out1),
	.prn(vcc));
defparam altera_reset_synchronizer_int_chain_out.is_wysiwyg = "true";
defparam altera_reset_synchronizer_int_chain_out.power_up = "low";

cyclonev_lcell_comb \altera_reset_synchronizer_int_chain[1]~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(altera_reset_synchronizer_int_chain_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \altera_reset_synchronizer_int_chain[1]~0 .extended_lut = "off";
defparam \altera_reset_synchronizer_int_chain[1]~0 .lut_mask = 64'h0000000000000000;
defparam \altera_reset_synchronizer_int_chain[1]~0 .shared_arith = "off";

dffeas \altera_reset_synchronizer_int_chain[1] (
	.clk(clk),
	.d(altera_reset_synchronizer_int_chain_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[1]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[1] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[1] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[0] (
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[0]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[0] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[0] .power_up = "low";

endmodule

module first_nios2_system_altera_reset_synchronizer_1 (
	altera_reset_synchronizer_int_chain_out1,
	clk,
	reset_reset_n)/* synthesis synthesis_greybox=1 */;
output 	altera_reset_synchronizer_int_chain_out1;
input 	clk;
input 	reset_reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \altera_reset_synchronizer_int_chain[1]~q ;
wire \altera_reset_synchronizer_int_chain[0]~q ;


dffeas altera_reset_synchronizer_int_chain_out(
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[0]~q ),
	.asdata(vcc),
	.clrn(reset_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(altera_reset_synchronizer_int_chain_out1),
	.prn(vcc));
defparam altera_reset_synchronizer_int_chain_out.is_wysiwyg = "true";
defparam altera_reset_synchronizer_int_chain_out.power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[1] (
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(reset_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[1]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[1] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[1] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[0] (
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[1]~q ),
	.asdata(vcc),
	.clrn(reset_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[0]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[0] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[0] .power_up = "low";

endmodule

module first_nios2_system_first_nios2_system_camData1 (
	readdata_0,
	readdata_1,
	readdata_2,
	readdata_3,
	readdata_4,
	readdata_5,
	readdata_6,
	A_mem_baddr_3,
	A_mem_baddr_2,
	Equal0,
	r_sync_rst,
	clk_clk,
	camdata1_external_connection_export_0,
	camdata1_external_connection_export_1,
	camdata1_external_connection_export_2,
	camdata1_external_connection_export_3,
	camdata1_external_connection_export_4,
	camdata1_external_connection_export_5,
	camdata1_external_connection_export_6)/* synthesis synthesis_greybox=1 */;
output 	readdata_0;
output 	readdata_1;
output 	readdata_2;
output 	readdata_3;
output 	readdata_4;
output 	readdata_5;
output 	readdata_6;
input 	A_mem_baddr_3;
input 	A_mem_baddr_2;
output 	Equal0;
input 	r_sync_rst;
input 	clk_clk;
input 	camdata1_external_connection_export_0;
input 	camdata1_external_connection_export_1;
input 	camdata1_external_connection_export_2;
input 	camdata1_external_connection_export_3;
input 	camdata1_external_connection_export_4;
input 	camdata1_external_connection_export_5;
input 	camdata1_external_connection_export_6;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \readdata[0] (
	.clk(clk_clk),
	.d(camdata1_external_connection_export_0),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(Equal0),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_0),
	.prn(vcc));
defparam \readdata[0] .is_wysiwyg = "true";
defparam \readdata[0] .power_up = "low";

dffeas \readdata[1] (
	.clk(clk_clk),
	.d(camdata1_external_connection_export_1),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(Equal0),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_1),
	.prn(vcc));
defparam \readdata[1] .is_wysiwyg = "true";
defparam \readdata[1] .power_up = "low";

dffeas \readdata[2] (
	.clk(clk_clk),
	.d(camdata1_external_connection_export_2),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(Equal0),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_2),
	.prn(vcc));
defparam \readdata[2] .is_wysiwyg = "true";
defparam \readdata[2] .power_up = "low";

dffeas \readdata[3] (
	.clk(clk_clk),
	.d(camdata1_external_connection_export_3),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(Equal0),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_3),
	.prn(vcc));
defparam \readdata[3] .is_wysiwyg = "true";
defparam \readdata[3] .power_up = "low";

dffeas \readdata[4] (
	.clk(clk_clk),
	.d(camdata1_external_connection_export_4),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(Equal0),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_4),
	.prn(vcc));
defparam \readdata[4] .is_wysiwyg = "true";
defparam \readdata[4] .power_up = "low";

dffeas \readdata[5] (
	.clk(clk_clk),
	.d(camdata1_external_connection_export_5),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(Equal0),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_5),
	.prn(vcc));
defparam \readdata[5] .is_wysiwyg = "true";
defparam \readdata[5] .power_up = "low";

dffeas \readdata[6] (
	.clk(clk_clk),
	.d(camdata1_external_connection_export_6),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(Equal0),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_6),
	.prn(vcc));
defparam \readdata[6] .is_wysiwyg = "true";
defparam \readdata[6] .power_up = "low";

cyclonev_lcell_comb \Equal0~0 (
	.dataa(!A_mem_baddr_3),
	.datab(!A_mem_baddr_2),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal0),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~0 .extended_lut = "off";
defparam \Equal0~0 .lut_mask = 64'h7777777777777777;
defparam \Equal0~0 .shared_arith = "off";

endmodule

module first_nios2_system_first_nios2_system_camData1_1 (
	readdata_0,
	readdata_1,
	readdata_2,
	readdata_3,
	readdata_4,
	readdata_5,
	readdata_6,
	Equal0,
	r_sync_rst,
	clk_clk,
	camdata2_external_connection_export_0,
	camdata2_external_connection_export_1,
	camdata2_external_connection_export_2,
	camdata2_external_connection_export_3,
	camdata2_external_connection_export_4,
	camdata2_external_connection_export_5,
	camdata2_external_connection_export_6)/* synthesis synthesis_greybox=1 */;
output 	readdata_0;
output 	readdata_1;
output 	readdata_2;
output 	readdata_3;
output 	readdata_4;
output 	readdata_5;
output 	readdata_6;
input 	Equal0;
input 	r_sync_rst;
input 	clk_clk;
input 	camdata2_external_connection_export_0;
input 	camdata2_external_connection_export_1;
input 	camdata2_external_connection_export_2;
input 	camdata2_external_connection_export_3;
input 	camdata2_external_connection_export_4;
input 	camdata2_external_connection_export_5;
input 	camdata2_external_connection_export_6;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \readdata[0] (
	.clk(clk_clk),
	.d(camdata2_external_connection_export_0),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(Equal0),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_0),
	.prn(vcc));
defparam \readdata[0] .is_wysiwyg = "true";
defparam \readdata[0] .power_up = "low";

dffeas \readdata[1] (
	.clk(clk_clk),
	.d(camdata2_external_connection_export_1),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(Equal0),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_1),
	.prn(vcc));
defparam \readdata[1] .is_wysiwyg = "true";
defparam \readdata[1] .power_up = "low";

dffeas \readdata[2] (
	.clk(clk_clk),
	.d(camdata2_external_connection_export_2),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(Equal0),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_2),
	.prn(vcc));
defparam \readdata[2] .is_wysiwyg = "true";
defparam \readdata[2] .power_up = "low";

dffeas \readdata[3] (
	.clk(clk_clk),
	.d(camdata2_external_connection_export_3),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(Equal0),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_3),
	.prn(vcc));
defparam \readdata[3] .is_wysiwyg = "true";
defparam \readdata[3] .power_up = "low";

dffeas \readdata[4] (
	.clk(clk_clk),
	.d(camdata2_external_connection_export_4),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(Equal0),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_4),
	.prn(vcc));
defparam \readdata[4] .is_wysiwyg = "true";
defparam \readdata[4] .power_up = "low";

dffeas \readdata[5] (
	.clk(clk_clk),
	.d(camdata2_external_connection_export_5),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(Equal0),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_5),
	.prn(vcc));
defparam \readdata[5] .is_wysiwyg = "true";
defparam \readdata[5] .power_up = "low";

dffeas \readdata[6] (
	.clk(clk_clk),
	.d(camdata2_external_connection_export_6),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(Equal0),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_6),
	.prn(vcc));
defparam \readdata[6] .is_wysiwyg = "true";
defparam \readdata[6] .power_up = "low";

endmodule

module first_nios2_system_first_nios2_system_camState1 (
	readdata_0,
	readdata_1,
	readdata_2,
	readdata_3,
	readdata_4,
	readdata_5,
	Equal0,
	r_sync_rst,
	clk_clk,
	camstate1_external_connection_export_0,
	camstate1_external_connection_export_1,
	camstate1_external_connection_export_2,
	camstate1_external_connection_export_3,
	camstate1_external_connection_export_4,
	camstate1_external_connection_export_5)/* synthesis synthesis_greybox=1 */;
output 	readdata_0;
output 	readdata_1;
output 	readdata_2;
output 	readdata_3;
output 	readdata_4;
output 	readdata_5;
input 	Equal0;
input 	r_sync_rst;
input 	clk_clk;
input 	camstate1_external_connection_export_0;
input 	camstate1_external_connection_export_1;
input 	camstate1_external_connection_export_2;
input 	camstate1_external_connection_export_3;
input 	camstate1_external_connection_export_4;
input 	camstate1_external_connection_export_5;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \readdata[0] (
	.clk(clk_clk),
	.d(camstate1_external_connection_export_0),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(Equal0),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_0),
	.prn(vcc));
defparam \readdata[0] .is_wysiwyg = "true";
defparam \readdata[0] .power_up = "low";

dffeas \readdata[1] (
	.clk(clk_clk),
	.d(camstate1_external_connection_export_1),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(Equal0),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_1),
	.prn(vcc));
defparam \readdata[1] .is_wysiwyg = "true";
defparam \readdata[1] .power_up = "low";

dffeas \readdata[2] (
	.clk(clk_clk),
	.d(camstate1_external_connection_export_2),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(Equal0),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_2),
	.prn(vcc));
defparam \readdata[2] .is_wysiwyg = "true";
defparam \readdata[2] .power_up = "low";

dffeas \readdata[3] (
	.clk(clk_clk),
	.d(camstate1_external_connection_export_3),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(Equal0),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_3),
	.prn(vcc));
defparam \readdata[3] .is_wysiwyg = "true";
defparam \readdata[3] .power_up = "low";

dffeas \readdata[4] (
	.clk(clk_clk),
	.d(camstate1_external_connection_export_4),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(Equal0),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_4),
	.prn(vcc));
defparam \readdata[4] .is_wysiwyg = "true";
defparam \readdata[4] .power_up = "low";

dffeas \readdata[5] (
	.clk(clk_clk),
	.d(camstate1_external_connection_export_5),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(Equal0),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_5),
	.prn(vcc));
defparam \readdata[5] .is_wysiwyg = "true";
defparam \readdata[5] .power_up = "low";

endmodule

module first_nios2_system_first_nios2_system_camState1_1 (
	readdata_0,
	readdata_1,
	readdata_2,
	readdata_3,
	readdata_4,
	readdata_5,
	Equal0,
	r_sync_rst,
	clk_clk,
	camstate2_external_connection_export_0,
	camstate2_external_connection_export_1,
	camstate2_external_connection_export_2,
	camstate2_external_connection_export_3,
	camstate2_external_connection_export_4,
	camstate2_external_connection_export_5)/* synthesis synthesis_greybox=1 */;
output 	readdata_0;
output 	readdata_1;
output 	readdata_2;
output 	readdata_3;
output 	readdata_4;
output 	readdata_5;
input 	Equal0;
input 	r_sync_rst;
input 	clk_clk;
input 	camstate2_external_connection_export_0;
input 	camstate2_external_connection_export_1;
input 	camstate2_external_connection_export_2;
input 	camstate2_external_connection_export_3;
input 	camstate2_external_connection_export_4;
input 	camstate2_external_connection_export_5;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \readdata[0] (
	.clk(clk_clk),
	.d(camstate2_external_connection_export_0),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(Equal0),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_0),
	.prn(vcc));
defparam \readdata[0] .is_wysiwyg = "true";
defparam \readdata[0] .power_up = "low";

dffeas \readdata[1] (
	.clk(clk_clk),
	.d(camstate2_external_connection_export_1),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(Equal0),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_1),
	.prn(vcc));
defparam \readdata[1] .is_wysiwyg = "true";
defparam \readdata[1] .power_up = "low";

dffeas \readdata[2] (
	.clk(clk_clk),
	.d(camstate2_external_connection_export_2),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(Equal0),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_2),
	.prn(vcc));
defparam \readdata[2] .is_wysiwyg = "true";
defparam \readdata[2] .power_up = "low";

dffeas \readdata[3] (
	.clk(clk_clk),
	.d(camstate2_external_connection_export_3),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(Equal0),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_3),
	.prn(vcc));
defparam \readdata[3] .is_wysiwyg = "true";
defparam \readdata[3] .power_up = "low";

dffeas \readdata[4] (
	.clk(clk_clk),
	.d(camstate2_external_connection_export_4),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(Equal0),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_4),
	.prn(vcc));
defparam \readdata[4] .is_wysiwyg = "true";
defparam \readdata[4] .power_up = "low";

dffeas \readdata[5] (
	.clk(clk_clk),
	.d(camstate2_external_connection_export_5),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(Equal0),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_5),
	.prn(vcc));
defparam \readdata[5] .is_wysiwyg = "true";
defparam \readdata[5] .power_up = "low";

endmodule

module first_nios2_system_first_nios2_system_cpu (
	av_readdata_pre_22,
	q_a_22,
	q_a_23,
	q_a_24,
	q_a_25,
	q_a_31,
	q_a_21,
	q_a_11,
	q_a_28,
	q_a_10,
	q_a_27,
	q_a_8,
	q_a_9,
	q_a_26,
	av_readdata_pre_20,
	q_a_20,
	av_readdata_pre_19,
	q_a_19,
	q_a_17,
	q_a_30,
	q_a_18,
	q_a_16,
	q_a_15,
	q_a_12,
	q_a_13,
	q_a_14,
	q_a_29,
	readdata_0,
	readdata_1,
	readdata_2,
	readdata_3,
	readdata_4,
	readdata_5,
	readdata_6,
	readdata_7,
	readdata_22,
	readdata_23,
	readdata_24,
	readdata_25,
	readdata_31,
	readdata_21,
	readdata_11,
	readdata_28,
	readdata_10,
	readdata_27,
	readdata_8,
	readdata_9,
	readdata_26,
	readdata_20,
	readdata_19,
	readdata_17,
	readdata_30,
	readdata_18,
	readdata_16,
	readdata_15,
	readdata_12,
	readdata_13,
	readdata_14,
	readdata_29,
	sr_0,
	ir_out_0,
	ir_out_1,
	A_st_data_0,
	A_mem_baddr_4,
	A_mem_baddr_5,
	A_mem_baddr_8,
	A_mem_baddr_16,
	A_mem_baddr_15,
	A_mem_baddr_14,
	A_mem_baddr_13,
	A_mem_baddr_12,
	A_mem_baddr_11,
	A_mem_baddr_10,
	A_mem_baddr_9,
	A_mem_baddr_7,
	A_mem_baddr_6,
	clr_break_line,
	d_write,
	A_mem_baddr_3,
	A_mem_baddr_2,
	r_sync_rst,
	A_st_data_1,
	A_st_data_2,
	A_st_data_3,
	A_st_data_4,
	A_st_data_5,
	A_st_data_6,
	A_st_data_7,
	d_read,
	W_debug_mode,
	read_latency_shift_reg_0,
	WideOr1,
	WideOr11,
	src0_valid,
	src0_valid1,
	read_latency_shift_reg_01,
	WideOr12,
	WideOr13,
	saved_grant_0,
	debug_mem_slave_waitrequest,
	mem_used_1,
	av_waitrequest,
	i_read,
	ic_fill_tag_5,
	ic_fill_tag_4,
	ic_fill_tag_3,
	ic_fill_tag_2,
	ic_fill_tag_1,
	ic_fill_tag_0,
	WideOr14,
	mem,
	timeout_occurred,
	control_register_0,
	av_readdata_9,
	av_readdata_8,
	src_payload,
	ic_fill_ap_offset_0,
	src_data_38,
	ic_fill_line_0,
	src_data_41,
	ic_fill_ap_offset_2,
	src_data_40,
	ic_fill_ap_offset_1,
	src_data_39,
	ic_fill_line_5,
	src_data_46,
	ic_fill_line_4,
	src_data_45,
	ic_fill_line_3,
	src_data_44,
	ic_fill_line_2,
	src_data_43,
	ic_fill_line_1,
	src_data_42,
	src_payload1,
	save_dest_id,
	WideOr0,
	nonposted_cmd_accepted,
	suppress_change_dest_id,
	r_early_rst,
	src_data_0,
	src_payload2,
	src_data_1,
	src_data_2,
	src_data_3,
	src_payload3,
	src_payload4,
	src_payload5,
	src_payload6,
	src_payload7,
	A_mem_byte_en_0,
	src_data_32,
	av_readdata_pre_221,
	src_payload8,
	av_readdata_pre_23,
	src_payload9,
	av_readdata_pre_24,
	src_payload10,
	av_readdata_pre_25,
	src_payload11,
	av_readdata_pre_31,
	src_payload12,
	av_readdata_pre_21,
	src_payload13,
	src_payload14,
	av_readdata_pre_11,
	src_payload15,
	src_payload16,
	av_readdata_pre_28,
	src_payload17,
	av_readdata_pre_10,
	src_payload18,
	src_payload19,
	av_readdata_pre_27,
	src_payload20,
	av_readdata_pre_8,
	src_payload21,
	src_payload22,
	av_readdata_pre_9,
	src_payload23,
	src_payload24,
	av_readdata_pre_26,
	src_payload25,
	av_readdata_pre_201,
	src_payload26,
	av_readdata_pre_191,
	src_payload27,
	av_readdata_pre_17,
	src_payload28,
	src_payload29,
	av_readdata_pre_30,
	src_payload30,
	av_readdata_pre_18,
	src_payload31,
	src_payload32,
	av_readdata_pre_16,
	src_payload33,
	src_payload34,
	av_readdata_pre_15,
	src_payload35,
	src_payload36,
	av_readdata_pre_12,
	src_payload37,
	src_payload38,
	av_readdata_pre_13,
	src_payload39,
	src_payload40,
	av_readdata_pre_14,
	src_payload41,
	src_payload42,
	av_readdata_pre_29,
	src_payload43,
	src_payload44,
	A_st_data_16,
	src_payload45,
	WideOr15,
	A_st_data_22,
	A_mem_byte_en_2,
	A_st_data_23,
	A_st_data_24,
	A_mem_byte_en_3,
	A_st_data_25,
	A_st_data_31,
	A_st_data_21,
	A_st_data_11,
	A_mem_byte_en_1,
	A_st_data_28,
	A_st_data_10,
	A_st_data_27,
	A_st_data_8,
	A_st_data_9,
	A_st_data_26,
	A_st_data_20,
	A_st_data_19,
	A_st_data_17,
	A_st_data_30,
	A_st_data_18,
	A_st_data_15,
	A_st_data_12,
	A_st_data_13,
	A_st_data_14,
	A_st_data_29,
	src_data_26,
	src_data_25,
	src_data_24,
	src_data_23,
	src_data_22,
	src_data_11,
	src_data_01,
	src_data_21,
	src_data_31,
	src_data_4,
	src_data_5,
	src_data_28,
	src_data_311,
	src_data_27,
	src_data_29,
	src_data_30,
	src_data_111,
	src_data_12,
	src_data_13,
	src_data_14,
	src_data_15,
	src_data_16,
	src_payload46,
	src_data_9,
	src_data_211,
	src_data_6,
	src_data_8,
	src_data_17,
	src_data_18,
	src_data_10,
	src_data_7,
	src_data_20,
	src_data_19,
	src_payload47,
	src_data_34,
	src_payload48,
	src_payload49,
	src_payload50,
	src_payload51,
	src_payload52,
	src_payload53,
	src_payload54,
	src_payload55,
	src_payload56,
	src_data_35,
	src_payload57,
	src_payload58,
	src_payload59,
	src_payload60,
	src_payload61,
	src_payload62,
	src_payload63,
	src_data_33,
	src_payload64,
	src_payload65,
	src_payload66,
	src_payload67,
	src_payload68,
	src_payload69,
	src_payload70,
	src_payload71,
	src_payload72,
	src_payload73,
	altera_internal_jtag,
	altera_internal_jtag1,
	state_1,
	state_4,
	virtual_ir_scan_reg,
	state_3,
	state_8,
	splitter_nodes_receive_1_3,
	irf_reg_0_2,
	irf_reg_1_2,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	av_readdata_pre_22;
input 	q_a_22;
input 	q_a_23;
input 	q_a_24;
input 	q_a_25;
input 	q_a_31;
input 	q_a_21;
input 	q_a_11;
input 	q_a_28;
input 	q_a_10;
input 	q_a_27;
input 	q_a_8;
input 	q_a_9;
input 	q_a_26;
input 	av_readdata_pre_20;
input 	q_a_20;
input 	av_readdata_pre_19;
input 	q_a_19;
input 	q_a_17;
input 	q_a_30;
input 	q_a_18;
input 	q_a_16;
input 	q_a_15;
input 	q_a_12;
input 	q_a_13;
input 	q_a_14;
input 	q_a_29;
output 	readdata_0;
output 	readdata_1;
output 	readdata_2;
output 	readdata_3;
output 	readdata_4;
output 	readdata_5;
output 	readdata_6;
output 	readdata_7;
output 	readdata_22;
output 	readdata_23;
output 	readdata_24;
output 	readdata_25;
output 	readdata_31;
output 	readdata_21;
output 	readdata_11;
output 	readdata_28;
output 	readdata_10;
output 	readdata_27;
output 	readdata_8;
output 	readdata_9;
output 	readdata_26;
output 	readdata_20;
output 	readdata_19;
output 	readdata_17;
output 	readdata_30;
output 	readdata_18;
output 	readdata_16;
output 	readdata_15;
output 	readdata_12;
output 	readdata_13;
output 	readdata_14;
output 	readdata_29;
output 	sr_0;
output 	ir_out_0;
output 	ir_out_1;
output 	A_st_data_0;
output 	A_mem_baddr_4;
output 	A_mem_baddr_5;
output 	A_mem_baddr_8;
output 	A_mem_baddr_16;
output 	A_mem_baddr_15;
output 	A_mem_baddr_14;
output 	A_mem_baddr_13;
output 	A_mem_baddr_12;
output 	A_mem_baddr_11;
output 	A_mem_baddr_10;
output 	A_mem_baddr_9;
output 	A_mem_baddr_7;
output 	A_mem_baddr_6;
output 	clr_break_line;
output 	d_write;
output 	A_mem_baddr_3;
output 	A_mem_baddr_2;
input 	r_sync_rst;
output 	A_st_data_1;
output 	A_st_data_2;
output 	A_st_data_3;
output 	A_st_data_4;
output 	A_st_data_5;
output 	A_st_data_6;
output 	A_st_data_7;
output 	d_read;
output 	W_debug_mode;
input 	read_latency_shift_reg_0;
input 	WideOr1;
input 	WideOr11;
input 	src0_valid;
input 	src0_valid1;
input 	read_latency_shift_reg_01;
input 	WideOr12;
input 	WideOr13;
input 	saved_grant_0;
output 	debug_mem_slave_waitrequest;
input 	mem_used_1;
input 	av_waitrequest;
output 	i_read;
output 	ic_fill_tag_5;
output 	ic_fill_tag_4;
output 	ic_fill_tag_3;
output 	ic_fill_tag_2;
output 	ic_fill_tag_1;
output 	ic_fill_tag_0;
input 	WideOr14;
input 	mem;
input 	timeout_occurred;
input 	control_register_0;
input 	av_readdata_9;
input 	av_readdata_8;
input 	src_payload;
output 	ic_fill_ap_offset_0;
input 	src_data_38;
output 	ic_fill_line_0;
input 	src_data_41;
output 	ic_fill_ap_offset_2;
input 	src_data_40;
output 	ic_fill_ap_offset_1;
input 	src_data_39;
output 	ic_fill_line_5;
input 	src_data_46;
output 	ic_fill_line_4;
input 	src_data_45;
output 	ic_fill_line_3;
input 	src_data_44;
output 	ic_fill_line_2;
input 	src_data_43;
output 	ic_fill_line_1;
input 	src_data_42;
input 	src_payload1;
input 	save_dest_id;
input 	WideOr0;
input 	nonposted_cmd_accepted;
input 	suppress_change_dest_id;
input 	r_early_rst;
input 	src_data_0;
input 	src_payload2;
input 	src_data_1;
input 	src_data_2;
input 	src_data_3;
input 	src_payload3;
input 	src_payload4;
input 	src_payload5;
input 	src_payload6;
input 	src_payload7;
output 	A_mem_byte_en_0;
input 	src_data_32;
input 	av_readdata_pre_221;
input 	src_payload8;
input 	av_readdata_pre_23;
input 	src_payload9;
input 	av_readdata_pre_24;
input 	src_payload10;
input 	av_readdata_pre_25;
input 	src_payload11;
input 	av_readdata_pre_31;
input 	src_payload12;
input 	av_readdata_pre_21;
input 	src_payload13;
input 	src_payload14;
input 	av_readdata_pre_11;
input 	src_payload15;
input 	src_payload16;
input 	av_readdata_pre_28;
input 	src_payload17;
input 	av_readdata_pre_10;
input 	src_payload18;
input 	src_payload19;
input 	av_readdata_pre_27;
input 	src_payload20;
input 	av_readdata_pre_8;
input 	src_payload21;
input 	src_payload22;
input 	av_readdata_pre_9;
input 	src_payload23;
input 	src_payload24;
input 	av_readdata_pre_26;
input 	src_payload25;
input 	av_readdata_pre_201;
input 	src_payload26;
input 	av_readdata_pre_191;
input 	src_payload27;
input 	av_readdata_pre_17;
input 	src_payload28;
input 	src_payload29;
input 	av_readdata_pre_30;
input 	src_payload30;
input 	av_readdata_pre_18;
input 	src_payload31;
input 	src_payload32;
input 	av_readdata_pre_16;
input 	src_payload33;
input 	src_payload34;
input 	av_readdata_pre_15;
input 	src_payload35;
input 	src_payload36;
input 	av_readdata_pre_12;
input 	src_payload37;
input 	src_payload38;
input 	av_readdata_pre_13;
input 	src_payload39;
input 	src_payload40;
input 	av_readdata_pre_14;
input 	src_payload41;
input 	src_payload42;
input 	av_readdata_pre_29;
input 	src_payload43;
input 	src_payload44;
output 	A_st_data_16;
input 	src_payload45;
input 	WideOr15;
output 	A_st_data_22;
output 	A_mem_byte_en_2;
output 	A_st_data_23;
output 	A_st_data_24;
output 	A_mem_byte_en_3;
output 	A_st_data_25;
output 	A_st_data_31;
output 	A_st_data_21;
output 	A_st_data_11;
output 	A_mem_byte_en_1;
output 	A_st_data_28;
output 	A_st_data_10;
output 	A_st_data_27;
output 	A_st_data_8;
output 	A_st_data_9;
output 	A_st_data_26;
output 	A_st_data_20;
output 	A_st_data_19;
output 	A_st_data_17;
output 	A_st_data_30;
output 	A_st_data_18;
output 	A_st_data_15;
output 	A_st_data_12;
output 	A_st_data_13;
output 	A_st_data_14;
output 	A_st_data_29;
input 	src_data_26;
input 	src_data_25;
input 	src_data_24;
input 	src_data_23;
input 	src_data_22;
input 	src_data_11;
input 	src_data_01;
input 	src_data_21;
input 	src_data_31;
input 	src_data_4;
input 	src_data_5;
input 	src_data_28;
input 	src_data_311;
input 	src_data_27;
input 	src_data_29;
input 	src_data_30;
input 	src_data_111;
input 	src_data_12;
input 	src_data_13;
input 	src_data_14;
input 	src_data_15;
input 	src_data_16;
input 	src_payload46;
input 	src_data_9;
input 	src_data_211;
input 	src_data_6;
input 	src_data_8;
input 	src_data_17;
input 	src_data_18;
input 	src_data_10;
input 	src_data_7;
input 	src_data_20;
input 	src_data_19;
input 	src_payload47;
input 	src_data_34;
input 	src_payload48;
input 	src_payload49;
input 	src_payload50;
input 	src_payload51;
input 	src_payload52;
input 	src_payload53;
input 	src_payload54;
input 	src_payload55;
input 	src_payload56;
input 	src_data_35;
input 	src_payload57;
input 	src_payload58;
input 	src_payload59;
input 	src_payload60;
input 	src_payload61;
input 	src_payload62;
input 	src_payload63;
input 	src_data_33;
input 	src_payload64;
input 	src_payload65;
input 	src_payload66;
input 	src_payload67;
input 	src_payload68;
input 	src_payload69;
input 	src_payload70;
input 	src_payload71;
input 	src_payload72;
input 	src_payload73;
input 	altera_internal_jtag;
input 	altera_internal_jtag1;
input 	state_1;
input 	state_4;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_8;
input 	splitter_nodes_receive_1_3;
input 	irf_reg_0_2;
input 	irf_reg_1_2;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



first_nios2_system_first_nios2_system_cpu_cpu cpu(
	.av_readdata_pre_22(av_readdata_pre_22),
	.q_a_22(q_a_22),
	.q_a_23(q_a_23),
	.q_a_24(q_a_24),
	.q_a_25(q_a_25),
	.q_a_31(q_a_31),
	.q_a_21(q_a_21),
	.q_a_11(q_a_11),
	.q_a_28(q_a_28),
	.q_a_10(q_a_10),
	.q_a_27(q_a_27),
	.q_a_8(q_a_8),
	.q_a_9(q_a_9),
	.q_a_26(q_a_26),
	.av_readdata_pre_20(av_readdata_pre_20),
	.q_a_20(q_a_20),
	.av_readdata_pre_19(av_readdata_pre_19),
	.q_a_19(q_a_19),
	.q_a_17(q_a_17),
	.q_a_30(q_a_30),
	.q_a_18(q_a_18),
	.q_a_16(q_a_16),
	.q_a_15(q_a_15),
	.q_a_12(q_a_12),
	.q_a_13(q_a_13),
	.q_a_14(q_a_14),
	.q_a_29(q_a_29),
	.readdata_0(readdata_0),
	.readdata_1(readdata_1),
	.readdata_2(readdata_2),
	.readdata_3(readdata_3),
	.readdata_4(readdata_4),
	.readdata_5(readdata_5),
	.readdata_6(readdata_6),
	.readdata_7(readdata_7),
	.readdata_22(readdata_22),
	.readdata_23(readdata_23),
	.readdata_24(readdata_24),
	.readdata_25(readdata_25),
	.readdata_31(readdata_31),
	.readdata_21(readdata_21),
	.readdata_11(readdata_11),
	.readdata_28(readdata_28),
	.readdata_10(readdata_10),
	.readdata_27(readdata_27),
	.readdata_8(readdata_8),
	.readdata_9(readdata_9),
	.readdata_26(readdata_26),
	.readdata_20(readdata_20),
	.readdata_19(readdata_19),
	.readdata_17(readdata_17),
	.readdata_30(readdata_30),
	.readdata_18(readdata_18),
	.readdata_16(readdata_16),
	.readdata_15(readdata_15),
	.readdata_12(readdata_12),
	.readdata_13(readdata_13),
	.readdata_14(readdata_14),
	.readdata_29(readdata_29),
	.sr_0(sr_0),
	.ir_out_0(ir_out_0),
	.ir_out_1(ir_out_1),
	.A_st_data_0(A_st_data_0),
	.A_mem_baddr_4(A_mem_baddr_4),
	.A_mem_baddr_5(A_mem_baddr_5),
	.A_mem_baddr_8(A_mem_baddr_8),
	.A_mem_baddr_16(A_mem_baddr_16),
	.A_mem_baddr_15(A_mem_baddr_15),
	.A_mem_baddr_14(A_mem_baddr_14),
	.A_mem_baddr_13(A_mem_baddr_13),
	.A_mem_baddr_12(A_mem_baddr_12),
	.A_mem_baddr_11(A_mem_baddr_11),
	.A_mem_baddr_10(A_mem_baddr_10),
	.A_mem_baddr_9(A_mem_baddr_9),
	.A_mem_baddr_7(A_mem_baddr_7),
	.A_mem_baddr_6(A_mem_baddr_6),
	.clr_break_line1(clr_break_line),
	.d_write1(d_write),
	.A_mem_baddr_3(A_mem_baddr_3),
	.A_mem_baddr_2(A_mem_baddr_2),
	.r_sync_rst(r_sync_rst),
	.A_st_data_1(A_st_data_1),
	.A_st_data_2(A_st_data_2),
	.A_st_data_3(A_st_data_3),
	.A_st_data_4(A_st_data_4),
	.A_st_data_5(A_st_data_5),
	.A_st_data_6(A_st_data_6),
	.A_st_data_7(A_st_data_7),
	.d_read1(d_read),
	.W_debug_mode1(W_debug_mode),
	.read_latency_shift_reg_0(read_latency_shift_reg_0),
	.WideOr1(WideOr1),
	.WideOr11(WideOr11),
	.src0_valid(src0_valid),
	.src0_valid1(src0_valid1),
	.read_latency_shift_reg_01(read_latency_shift_reg_01),
	.WideOr12(WideOr12),
	.WideOr13(WideOr13),
	.saved_grant_0(saved_grant_0),
	.debug_mem_slave_waitrequest(debug_mem_slave_waitrequest),
	.mem_used_1(mem_used_1),
	.av_waitrequest(av_waitrequest),
	.i_read1(i_read),
	.ic_fill_tag_5(ic_fill_tag_5),
	.ic_fill_tag_4(ic_fill_tag_4),
	.ic_fill_tag_3(ic_fill_tag_3),
	.ic_fill_tag_2(ic_fill_tag_2),
	.ic_fill_tag_1(ic_fill_tag_1),
	.ic_fill_tag_0(ic_fill_tag_0),
	.WideOr14(WideOr14),
	.mem(mem),
	.timeout_occurred(timeout_occurred),
	.control_register_0(control_register_0),
	.av_readdata_9(av_readdata_9),
	.av_readdata_8(av_readdata_8),
	.src_payload(src_payload),
	.ic_fill_ap_offset_0(ic_fill_ap_offset_0),
	.src_data_38(src_data_38),
	.ic_fill_line_0(ic_fill_line_0),
	.src_data_41(src_data_41),
	.ic_fill_ap_offset_2(ic_fill_ap_offset_2),
	.src_data_40(src_data_40),
	.ic_fill_ap_offset_1(ic_fill_ap_offset_1),
	.src_data_39(src_data_39),
	.ic_fill_line_5(ic_fill_line_5),
	.src_data_46(src_data_46),
	.ic_fill_line_4(ic_fill_line_4),
	.src_data_45(src_data_45),
	.ic_fill_line_3(ic_fill_line_3),
	.src_data_44(src_data_44),
	.ic_fill_line_2(ic_fill_line_2),
	.src_data_43(src_data_43),
	.ic_fill_line_1(ic_fill_line_1),
	.src_data_42(src_data_42),
	.src_payload1(src_payload1),
	.save_dest_id(save_dest_id),
	.WideOr0(WideOr0),
	.nonposted_cmd_accepted(nonposted_cmd_accepted),
	.suppress_change_dest_id(suppress_change_dest_id),
	.r_early_rst(r_early_rst),
	.d_readdata({src_payload12,src_payload30,src_payload43,src_payload17,src_payload20,src_payload25,src_payload11,src_payload10,src_payload9,src_payload8,src_payload14,src_payload26,src_payload27,src_payload32,src_payload29,src_payload34,src_payload36,src_payload42,src_payload40,
src_payload38,src_payload16,src_payload19,src_payload24,src_payload22,src_payload6,src_payload5,src_payload4,src_payload3,src_data_3,src_data_2,src_data_1,src_data_0}),
	.src_payload2(src_payload2),
	.src_payload3(src_payload7),
	.A_mem_byte_en_0(A_mem_byte_en_0),
	.src_data_32(src_data_32),
	.av_readdata_pre_221(av_readdata_pre_221),
	.av_readdata_pre_23(av_readdata_pre_23),
	.av_readdata_pre_24(av_readdata_pre_24),
	.av_readdata_pre_25(av_readdata_pre_25),
	.av_readdata_pre_31(av_readdata_pre_31),
	.av_readdata_pre_21(av_readdata_pre_21),
	.src_payload4(src_payload13),
	.av_readdata_pre_11(av_readdata_pre_11),
	.src_payload5(src_payload15),
	.av_readdata_pre_28(av_readdata_pre_28),
	.av_readdata_pre_10(av_readdata_pre_10),
	.src_payload6(src_payload18),
	.av_readdata_pre_27(av_readdata_pre_27),
	.av_readdata_pre_8(av_readdata_pre_8),
	.src_payload7(src_payload21),
	.av_readdata_pre_9(av_readdata_pre_9),
	.src_payload8(src_payload23),
	.av_readdata_pre_26(av_readdata_pre_26),
	.av_readdata_pre_201(av_readdata_pre_201),
	.av_readdata_pre_191(av_readdata_pre_191),
	.av_readdata_pre_17(av_readdata_pre_17),
	.src_payload9(src_payload28),
	.av_readdata_pre_30(av_readdata_pre_30),
	.av_readdata_pre_18(av_readdata_pre_18),
	.src_payload10(src_payload31),
	.av_readdata_pre_16(av_readdata_pre_16),
	.src_payload11(src_payload33),
	.av_readdata_pre_15(av_readdata_pre_15),
	.src_payload12(src_payload35),
	.av_readdata_pre_12(av_readdata_pre_12),
	.src_payload13(src_payload37),
	.av_readdata_pre_13(av_readdata_pre_13),
	.src_payload14(src_payload39),
	.av_readdata_pre_14(av_readdata_pre_14),
	.src_payload15(src_payload41),
	.av_readdata_pre_29(av_readdata_pre_29),
	.src_payload16(src_payload44),
	.A_st_data_16(A_st_data_16),
	.src_payload17(src_payload45),
	.WideOr15(WideOr15),
	.A_st_data_22(A_st_data_22),
	.A_mem_byte_en_2(A_mem_byte_en_2),
	.A_st_data_23(A_st_data_23),
	.A_st_data_24(A_st_data_24),
	.A_mem_byte_en_3(A_mem_byte_en_3),
	.A_st_data_25(A_st_data_25),
	.A_st_data_31(A_st_data_31),
	.A_st_data_21(A_st_data_21),
	.A_st_data_11(A_st_data_11),
	.A_mem_byte_en_1(A_mem_byte_en_1),
	.A_st_data_28(A_st_data_28),
	.A_st_data_10(A_st_data_10),
	.A_st_data_27(A_st_data_27),
	.A_st_data_8(A_st_data_8),
	.A_st_data_9(A_st_data_9),
	.A_st_data_26(A_st_data_26),
	.A_st_data_20(A_st_data_20),
	.A_st_data_19(A_st_data_19),
	.A_st_data_17(A_st_data_17),
	.A_st_data_30(A_st_data_30),
	.A_st_data_18(A_st_data_18),
	.A_st_data_15(A_st_data_15),
	.A_st_data_12(A_st_data_12),
	.A_st_data_13(A_st_data_13),
	.A_st_data_14(A_st_data_14),
	.A_st_data_29(A_st_data_29),
	.i_readdata({src_data_311,src_data_30,src_data_29,src_data_28,src_data_27,src_data_26,src_data_25,src_data_24,src_data_23,src_data_22,src_data_211,src_data_20,src_data_19,src_data_18,src_data_17,src_data_16,src_data_15,src_data_14,src_data_13,src_data_12,src_data_111,src_data_10,src_data_9,
src_data_8,src_data_7,src_data_6,src_data_5,src_data_4,src_data_31,src_data_21,src_data_11,src_data_01}),
	.src_payload18(src_payload46),
	.src_payload19(src_payload47),
	.src_data_34(src_data_34),
	.src_payload20(src_payload48),
	.src_payload21(src_payload49),
	.src_payload22(src_payload50),
	.src_payload23(src_payload51),
	.src_payload24(src_payload52),
	.src_payload25(src_payload53),
	.src_payload26(src_payload54),
	.src_payload27(src_payload55),
	.src_payload28(src_payload56),
	.src_data_35(src_data_35),
	.src_payload29(src_payload57),
	.src_payload30(src_payload58),
	.src_payload31(src_payload59),
	.src_payload32(src_payload60),
	.src_payload33(src_payload61),
	.src_payload34(src_payload62),
	.src_payload35(src_payload63),
	.src_data_33(src_data_33),
	.src_payload36(src_payload64),
	.src_payload37(src_payload65),
	.src_payload38(src_payload66),
	.src_payload39(src_payload67),
	.src_payload40(src_payload68),
	.src_payload41(src_payload69),
	.src_payload42(src_payload70),
	.src_payload43(src_payload71),
	.src_payload44(src_payload72),
	.src_payload45(src_payload73),
	.altera_internal_jtag(altera_internal_jtag),
	.altera_internal_jtag1(altera_internal_jtag1),
	.state_1(state_1),
	.state_4(state_4),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.state_8(state_8),
	.splitter_nodes_receive_1_3(splitter_nodes_receive_1_3),
	.irf_reg_0_2(irf_reg_0_2),
	.irf_reg_1_2(irf_reg_1_2),
	.clk_clk(clk_clk));

endmodule

module first_nios2_system_first_nios2_system_cpu_cpu (
	av_readdata_pre_22,
	q_a_22,
	q_a_23,
	q_a_24,
	q_a_25,
	q_a_31,
	q_a_21,
	q_a_11,
	q_a_28,
	q_a_10,
	q_a_27,
	q_a_8,
	q_a_9,
	q_a_26,
	av_readdata_pre_20,
	q_a_20,
	av_readdata_pre_19,
	q_a_19,
	q_a_17,
	q_a_30,
	q_a_18,
	q_a_16,
	q_a_15,
	q_a_12,
	q_a_13,
	q_a_14,
	q_a_29,
	readdata_0,
	readdata_1,
	readdata_2,
	readdata_3,
	readdata_4,
	readdata_5,
	readdata_6,
	readdata_7,
	readdata_22,
	readdata_23,
	readdata_24,
	readdata_25,
	readdata_31,
	readdata_21,
	readdata_11,
	readdata_28,
	readdata_10,
	readdata_27,
	readdata_8,
	readdata_9,
	readdata_26,
	readdata_20,
	readdata_19,
	readdata_17,
	readdata_30,
	readdata_18,
	readdata_16,
	readdata_15,
	readdata_12,
	readdata_13,
	readdata_14,
	readdata_29,
	sr_0,
	ir_out_0,
	ir_out_1,
	A_st_data_0,
	A_mem_baddr_4,
	A_mem_baddr_5,
	A_mem_baddr_8,
	A_mem_baddr_16,
	A_mem_baddr_15,
	A_mem_baddr_14,
	A_mem_baddr_13,
	A_mem_baddr_12,
	A_mem_baddr_11,
	A_mem_baddr_10,
	A_mem_baddr_9,
	A_mem_baddr_7,
	A_mem_baddr_6,
	clr_break_line1,
	d_write1,
	A_mem_baddr_3,
	A_mem_baddr_2,
	r_sync_rst,
	A_st_data_1,
	A_st_data_2,
	A_st_data_3,
	A_st_data_4,
	A_st_data_5,
	A_st_data_6,
	A_st_data_7,
	d_read1,
	W_debug_mode1,
	read_latency_shift_reg_0,
	WideOr1,
	WideOr11,
	src0_valid,
	src0_valid1,
	read_latency_shift_reg_01,
	WideOr12,
	WideOr13,
	saved_grant_0,
	debug_mem_slave_waitrequest,
	mem_used_1,
	av_waitrequest,
	i_read1,
	ic_fill_tag_5,
	ic_fill_tag_4,
	ic_fill_tag_3,
	ic_fill_tag_2,
	ic_fill_tag_1,
	ic_fill_tag_0,
	WideOr14,
	mem,
	timeout_occurred,
	control_register_0,
	av_readdata_9,
	av_readdata_8,
	src_payload,
	ic_fill_ap_offset_0,
	src_data_38,
	ic_fill_line_0,
	src_data_41,
	ic_fill_ap_offset_2,
	src_data_40,
	ic_fill_ap_offset_1,
	src_data_39,
	ic_fill_line_5,
	src_data_46,
	ic_fill_line_4,
	src_data_45,
	ic_fill_line_3,
	src_data_44,
	ic_fill_line_2,
	src_data_43,
	ic_fill_line_1,
	src_data_42,
	src_payload1,
	save_dest_id,
	WideOr0,
	nonposted_cmd_accepted,
	suppress_change_dest_id,
	r_early_rst,
	d_readdata,
	src_payload2,
	src_payload3,
	A_mem_byte_en_0,
	src_data_32,
	av_readdata_pre_221,
	av_readdata_pre_23,
	av_readdata_pre_24,
	av_readdata_pre_25,
	av_readdata_pre_31,
	av_readdata_pre_21,
	src_payload4,
	av_readdata_pre_11,
	src_payload5,
	av_readdata_pre_28,
	av_readdata_pre_10,
	src_payload6,
	av_readdata_pre_27,
	av_readdata_pre_8,
	src_payload7,
	av_readdata_pre_9,
	src_payload8,
	av_readdata_pre_26,
	av_readdata_pre_201,
	av_readdata_pre_191,
	av_readdata_pre_17,
	src_payload9,
	av_readdata_pre_30,
	av_readdata_pre_18,
	src_payload10,
	av_readdata_pre_16,
	src_payload11,
	av_readdata_pre_15,
	src_payload12,
	av_readdata_pre_12,
	src_payload13,
	av_readdata_pre_13,
	src_payload14,
	av_readdata_pre_14,
	src_payload15,
	av_readdata_pre_29,
	src_payload16,
	A_st_data_16,
	src_payload17,
	WideOr15,
	A_st_data_22,
	A_mem_byte_en_2,
	A_st_data_23,
	A_st_data_24,
	A_mem_byte_en_3,
	A_st_data_25,
	A_st_data_31,
	A_st_data_21,
	A_st_data_11,
	A_mem_byte_en_1,
	A_st_data_28,
	A_st_data_10,
	A_st_data_27,
	A_st_data_8,
	A_st_data_9,
	A_st_data_26,
	A_st_data_20,
	A_st_data_19,
	A_st_data_17,
	A_st_data_30,
	A_st_data_18,
	A_st_data_15,
	A_st_data_12,
	A_st_data_13,
	A_st_data_14,
	A_st_data_29,
	i_readdata,
	src_payload18,
	src_payload19,
	src_data_34,
	src_payload20,
	src_payload21,
	src_payload22,
	src_payload23,
	src_payload24,
	src_payload25,
	src_payload26,
	src_payload27,
	src_payload28,
	src_data_35,
	src_payload29,
	src_payload30,
	src_payload31,
	src_payload32,
	src_payload33,
	src_payload34,
	src_payload35,
	src_data_33,
	src_payload36,
	src_payload37,
	src_payload38,
	src_payload39,
	src_payload40,
	src_payload41,
	src_payload42,
	src_payload43,
	src_payload44,
	src_payload45,
	altera_internal_jtag,
	altera_internal_jtag1,
	state_1,
	state_4,
	virtual_ir_scan_reg,
	state_3,
	state_8,
	splitter_nodes_receive_1_3,
	irf_reg_0_2,
	irf_reg_1_2,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	av_readdata_pre_22;
input 	q_a_22;
input 	q_a_23;
input 	q_a_24;
input 	q_a_25;
input 	q_a_31;
input 	q_a_21;
input 	q_a_11;
input 	q_a_28;
input 	q_a_10;
input 	q_a_27;
input 	q_a_8;
input 	q_a_9;
input 	q_a_26;
input 	av_readdata_pre_20;
input 	q_a_20;
input 	av_readdata_pre_19;
input 	q_a_19;
input 	q_a_17;
input 	q_a_30;
input 	q_a_18;
input 	q_a_16;
input 	q_a_15;
input 	q_a_12;
input 	q_a_13;
input 	q_a_14;
input 	q_a_29;
output 	readdata_0;
output 	readdata_1;
output 	readdata_2;
output 	readdata_3;
output 	readdata_4;
output 	readdata_5;
output 	readdata_6;
output 	readdata_7;
output 	readdata_22;
output 	readdata_23;
output 	readdata_24;
output 	readdata_25;
output 	readdata_31;
output 	readdata_21;
output 	readdata_11;
output 	readdata_28;
output 	readdata_10;
output 	readdata_27;
output 	readdata_8;
output 	readdata_9;
output 	readdata_26;
output 	readdata_20;
output 	readdata_19;
output 	readdata_17;
output 	readdata_30;
output 	readdata_18;
output 	readdata_16;
output 	readdata_15;
output 	readdata_12;
output 	readdata_13;
output 	readdata_14;
output 	readdata_29;
output 	sr_0;
output 	ir_out_0;
output 	ir_out_1;
output 	A_st_data_0;
output 	A_mem_baddr_4;
output 	A_mem_baddr_5;
output 	A_mem_baddr_8;
output 	A_mem_baddr_16;
output 	A_mem_baddr_15;
output 	A_mem_baddr_14;
output 	A_mem_baddr_13;
output 	A_mem_baddr_12;
output 	A_mem_baddr_11;
output 	A_mem_baddr_10;
output 	A_mem_baddr_9;
output 	A_mem_baddr_7;
output 	A_mem_baddr_6;
output 	clr_break_line1;
output 	d_write1;
output 	A_mem_baddr_3;
output 	A_mem_baddr_2;
input 	r_sync_rst;
output 	A_st_data_1;
output 	A_st_data_2;
output 	A_st_data_3;
output 	A_st_data_4;
output 	A_st_data_5;
output 	A_st_data_6;
output 	A_st_data_7;
output 	d_read1;
output 	W_debug_mode1;
input 	read_latency_shift_reg_0;
input 	WideOr1;
input 	WideOr11;
input 	src0_valid;
input 	src0_valid1;
input 	read_latency_shift_reg_01;
input 	WideOr12;
input 	WideOr13;
input 	saved_grant_0;
output 	debug_mem_slave_waitrequest;
input 	mem_used_1;
input 	av_waitrequest;
output 	i_read1;
output 	ic_fill_tag_5;
output 	ic_fill_tag_4;
output 	ic_fill_tag_3;
output 	ic_fill_tag_2;
output 	ic_fill_tag_1;
output 	ic_fill_tag_0;
input 	WideOr14;
input 	mem;
input 	timeout_occurred;
input 	control_register_0;
input 	av_readdata_9;
input 	av_readdata_8;
input 	src_payload;
output 	ic_fill_ap_offset_0;
input 	src_data_38;
output 	ic_fill_line_0;
input 	src_data_41;
output 	ic_fill_ap_offset_2;
input 	src_data_40;
output 	ic_fill_ap_offset_1;
input 	src_data_39;
output 	ic_fill_line_5;
input 	src_data_46;
output 	ic_fill_line_4;
input 	src_data_45;
output 	ic_fill_line_3;
input 	src_data_44;
output 	ic_fill_line_2;
input 	src_data_43;
output 	ic_fill_line_1;
input 	src_data_42;
input 	src_payload1;
input 	save_dest_id;
input 	WideOr0;
input 	nonposted_cmd_accepted;
input 	suppress_change_dest_id;
input 	r_early_rst;
input 	[31:0] d_readdata;
input 	src_payload2;
input 	src_payload3;
output 	A_mem_byte_en_0;
input 	src_data_32;
input 	av_readdata_pre_221;
input 	av_readdata_pre_23;
input 	av_readdata_pre_24;
input 	av_readdata_pre_25;
input 	av_readdata_pre_31;
input 	av_readdata_pre_21;
input 	src_payload4;
input 	av_readdata_pre_11;
input 	src_payload5;
input 	av_readdata_pre_28;
input 	av_readdata_pre_10;
input 	src_payload6;
input 	av_readdata_pre_27;
input 	av_readdata_pre_8;
input 	src_payload7;
input 	av_readdata_pre_9;
input 	src_payload8;
input 	av_readdata_pre_26;
input 	av_readdata_pre_201;
input 	av_readdata_pre_191;
input 	av_readdata_pre_17;
input 	src_payload9;
input 	av_readdata_pre_30;
input 	av_readdata_pre_18;
input 	src_payload10;
input 	av_readdata_pre_16;
input 	src_payload11;
input 	av_readdata_pre_15;
input 	src_payload12;
input 	av_readdata_pre_12;
input 	src_payload13;
input 	av_readdata_pre_13;
input 	src_payload14;
input 	av_readdata_pre_14;
input 	src_payload15;
input 	av_readdata_pre_29;
input 	src_payload16;
output 	A_st_data_16;
input 	src_payload17;
input 	WideOr15;
output 	A_st_data_22;
output 	A_mem_byte_en_2;
output 	A_st_data_23;
output 	A_st_data_24;
output 	A_mem_byte_en_3;
output 	A_st_data_25;
output 	A_st_data_31;
output 	A_st_data_21;
output 	A_st_data_11;
output 	A_mem_byte_en_1;
output 	A_st_data_28;
output 	A_st_data_10;
output 	A_st_data_27;
output 	A_st_data_8;
output 	A_st_data_9;
output 	A_st_data_26;
output 	A_st_data_20;
output 	A_st_data_19;
output 	A_st_data_17;
output 	A_st_data_30;
output 	A_st_data_18;
output 	A_st_data_15;
output 	A_st_data_12;
output 	A_st_data_13;
output 	A_st_data_14;
output 	A_st_data_29;
input 	[31:0] i_readdata;
input 	src_payload18;
input 	src_payload19;
input 	src_data_34;
input 	src_payload20;
input 	src_payload21;
input 	src_payload22;
input 	src_payload23;
input 	src_payload24;
input 	src_payload25;
input 	src_payload26;
input 	src_payload27;
input 	src_payload28;
input 	src_data_35;
input 	src_payload29;
input 	src_payload30;
input 	src_payload31;
input 	src_payload32;
input 	src_payload33;
input 	src_payload34;
input 	src_payload35;
input 	src_data_33;
input 	src_payload36;
input 	src_payload37;
input 	src_payload38;
input 	src_payload39;
input 	src_payload40;
input 	src_payload41;
input 	src_payload42;
input 	src_payload43;
input 	src_payload44;
input 	src_payload45;
input 	altera_internal_jtag;
input 	altera_internal_jtag1;
input 	state_1;
input 	state_4;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_8;
input 	splitter_nodes_receive_1_3;
input 	irf_reg_0_2;
input 	irf_reg_1_2;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[0] ;
wire \first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[1] ;
wire \first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[2] ;
wire \first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[3] ;
wire \first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[4] ;
wire \first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[5] ;
wire \first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[6] ;
wire \first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[7] ;
wire \first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[3] ;
wire \first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[22] ;
wire \first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[22] ;
wire \first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[23] ;
wire \first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[23] ;
wire \first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[24] ;
wire \first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[24] ;
wire \first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[0] ;
wire \first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[25] ;
wire \first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[25] ;
wire \first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[2] ;
wire \first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[31] ;
wire \first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[31] ;
wire \first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[7] ;
wire \first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[21] ;
wire \first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[21] ;
wire \first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[11] ;
wire \first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[11] ;
wire \first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[28] ;
wire \first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[28] ;
wire \first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[10] ;
wire \first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[10] ;
wire \first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[27] ;
wire \first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[27] ;
wire \first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[8] ;
wire \first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[8] ;
wire \first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[9] ;
wire \first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[9] ;
wire \first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[4] ;
wire \first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[5] ;
wire \first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[6] ;
wire \first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[26] ;
wire \first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[26] ;
wire \first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[20] ;
wire \first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[20] ;
wire \first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[19] ;
wire \first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[19] ;
wire \first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[17] ;
wire \first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[17] ;
wire \first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[30] ;
wire \first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[30] ;
wire \first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[1] ;
wire \first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[18] ;
wire \first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[18] ;
wire \first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[16] ;
wire \first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[16] ;
wire \first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[15] ;
wire \first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[15] ;
wire \first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[12] ;
wire \first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[12] ;
wire \first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[13] ;
wire \first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[13] ;
wire \first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[14] ;
wire \first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[14] ;
wire \first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[29] ;
wire \first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[29] ;
wire \first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[26] ;
wire \first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[25] ;
wire \first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[24] ;
wire \first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[23] ;
wire \first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[22] ;
wire \first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[1] ;
wire \first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[0] ;
wire \first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[2] ;
wire \first_nios2_system_cpu_cpu_ic_tag|the_altsyncram|auto_generated|q_b[5] ;
wire \first_nios2_system_cpu_cpu_ic_tag|the_altsyncram|auto_generated|q_b[0] ;
wire \first_nios2_system_cpu_cpu_ic_tag|the_altsyncram|auto_generated|q_b[1] ;
wire \first_nios2_system_cpu_cpu_ic_tag|the_altsyncram|auto_generated|q_b[2] ;
wire \first_nios2_system_cpu_cpu_ic_tag|the_altsyncram|auto_generated|q_b[3] ;
wire \first_nios2_system_cpu_cpu_ic_tag|the_altsyncram|auto_generated|q_b[4] ;
wire \first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[3] ;
wire \first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[4] ;
wire \first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[5] ;
wire \first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[28] ;
wire \first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[31] ;
wire \first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[27] ;
wire \first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[29] ;
wire \first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[30] ;
wire \first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[11] ;
wire \first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[12] ;
wire \first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[13] ;
wire \first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[14] ;
wire \first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[15] ;
wire \first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[16] ;
wire \first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[9] ;
wire \first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[21] ;
wire \first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[6] ;
wire \first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[8] ;
wire \first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[17] ;
wire \first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[18] ;
wire \first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[10] ;
wire \first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[7] ;
wire \first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[20] ;
wire \first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[19] ;
wire \first_nios2_system_cpu_cpu_bht|the_altsyncram|auto_generated|q_b[1] ;
wire \first_nios2_system_cpu_cpu_ic_tag|the_altsyncram|auto_generated|q_b[11] ;
wire \first_nios2_system_cpu_cpu_ic_tag|the_altsyncram|auto_generated|q_b[13] ;
wire \first_nios2_system_cpu_cpu_ic_tag|the_altsyncram|auto_generated|q_b[10] ;
wire \first_nios2_system_cpu_cpu_ic_tag|the_altsyncram|auto_generated|q_b[12] ;
wire \ic_tag_wraddress[0]~q ;
wire \ic_tag_wraddress[1]~q ;
wire \ic_tag_wraddress[2]~q ;
wire \ic_tag_wraddress[3]~q ;
wire \ic_tag_wraddress[4]~q ;
wire \ic_tag_wraddress[5]~q ;
wire \ic_fill_valid_bits[5]~q ;
wire \ic_fill_valid_bits[7]~q ;
wire \ic_fill_valid_bits[4]~q ;
wire \first_nios2_system_cpu_cpu_ic_tag|the_altsyncram|auto_generated|q_b[7] ;
wire \first_nios2_system_cpu_cpu_ic_tag|the_altsyncram|auto_generated|q_b[9] ;
wire \first_nios2_system_cpu_cpu_ic_tag|the_altsyncram|auto_generated|q_b[6] ;
wire \first_nios2_system_cpu_cpu_ic_tag|the_altsyncram|auto_generated|q_b[8] ;
wire \ic_fill_valid_bits[6]~q ;
wire \ic_fill_valid_bits[1]~q ;
wire \ic_fill_valid_bits[3]~q ;
wire \ic_fill_valid_bits[0]~q ;
wire \ic_fill_valid_bits[2]~q ;
wire \first_nios2_system_cpu_cpu_bht|the_altsyncram|auto_generated|q_b[0] ;
wire \the_first_nios2_system_cpu_cpu_nios2_oci|the_first_nios2_system_cpu_cpu_nios2_avalon_reg|oci_single_step_mode~q ;
wire \the_first_nios2_system_cpu_cpu_nios2_oci|the_first_nios2_system_cpu_cpu_nios2_oci_debug|jtag_break~q ;
wire \the_first_nios2_system_cpu_cpu_nios2_oci|the_first_nios2_system_cpu_cpu_nios2_avalon_reg|oci_ienable[1]~q ;
wire \the_first_nios2_system_cpu_cpu_nios2_oci|the_first_nios2_system_cpu_cpu_nios2_avalon_reg|oci_ienable[16]~q ;
wire \rf_b_rd_port_addr[0]~0_combout ;
wire \rf_b_rd_port_addr[1]~1_combout ;
wire \rf_b_rd_port_addr[2]~2_combout ;
wire \rf_b_rd_port_addr[3]~3_combout ;
wire \rf_b_rd_port_addr[4]~4_combout ;
wire \the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[0]~q ;
wire \the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[1]~q ;
wire \the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[2]~q ;
wire \the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[3]~q ;
wire \the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[4]~q ;
wire \the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[5]~q ;
wire \the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[6]~q ;
wire \the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[7]~q ;
wire \rf_a_rd_port_addr[0]~0_combout ;
wire \rf_a_rd_port_addr[1]~1_combout ;
wire \rf_a_rd_port_addr[2]~2_combout ;
wire \rf_a_rd_port_addr[3]~3_combout ;
wire \rf_a_rd_port_addr[4]~4_combout ;
wire \the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[11]~q ;
wire \the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[10]~q ;
wire \the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[8]~q ;
wire \the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[9]~q ;
wire \the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[15]~q ;
wire \the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[12]~q ;
wire \the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[13]~q ;
wire \the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[14]~q ;
wire \i_readdata_d1[26]~q ;
wire \i_readdata_d1[25]~q ;
wire \i_readdata_d1[24]~q ;
wire \i_readdata_d1[23]~q ;
wire \i_readdata_d1[22]~q ;
wire \i_readdata_d1[1]~q ;
wire \i_readdata_d1[0]~q ;
wire \i_readdata_d1[2]~q ;
wire \ic_tag_clr_valid_bits~q ;
wire \ic_tag_wren~combout ;
wire \i_readdata_d1[3]~q ;
wire \i_readdata_d1[4]~q ;
wire \i_readdata_d1[5]~q ;
wire \i_readdata_d1[28]~q ;
wire \i_readdata_d1[31]~q ;
wire \i_readdata_d1[27]~q ;
wire \i_readdata_d1[29]~q ;
wire \i_readdata_d1[30]~q ;
wire \i_readdata_d1[11]~q ;
wire \i_readdata_d1[12]~q ;
wire \i_readdata_d1[13]~q ;
wire \i_readdata_d1[14]~q ;
wire \i_readdata_d1[15]~q ;
wire \i_readdata_d1[16]~q ;
wire \i_readdata_d1[9]~q ;
wire \the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p3|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[6]~q ;
wire \i_readdata_d1[21]~q ;
wire \the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p3|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[7]~q ;
wire \the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p3|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[8]~q ;
wire \i_readdata_d1[6]~q ;
wire \the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p3|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[9]~q ;
wire \i_readdata_d1[8]~q ;
wire \the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p3|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[15]~q ;
wire \the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p3|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[5]~q ;
wire \i_readdata_d1[17]~q ;
wire \the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p3|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[12]~q ;
wire \i_readdata_d1[18]~q ;
wire \the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p3|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[11]~q ;
wire \i_readdata_d1[10]~q ;
wire \the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p3|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[10]~q ;
wire \the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p3|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[4]~q ;
wire \the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p3|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[3]~q ;
wire \the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p3|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[1]~q ;
wire \i_readdata_d1[7]~q ;
wire \the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p3|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[14]~q ;
wire \i_readdata_d1[20]~q ;
wire \the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p3|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[2]~q ;
wire \the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p3|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[0]~q ;
wire \i_readdata_d1[19]~q ;
wire \the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p3|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[13]~q ;
wire \M_ctrl_br_cond~q ;
wire \M_bht_wr_en_unfiltered~combout ;
wire \M_bht_data[1]~q ;
wire \M_bht_data[0]~q ;
wire \M_br_mispredict~q ;
wire \M_bht_wr_data_unfiltered[1]~0_combout ;
wire \M_bht_ptr_unfiltered[0]~q ;
wire \M_bht_ptr_unfiltered[1]~q ;
wire \M_bht_ptr_unfiltered[2]~q ;
wire \M_bht_ptr_unfiltered[3]~q ;
wire \M_bht_ptr_unfiltered[4]~q ;
wire \M_bht_ptr_unfiltered[5]~q ;
wire \M_bht_ptr_unfiltered[6]~q ;
wire \M_bht_ptr_unfiltered[7]~q ;
wire \M_br_cond_taken_history[0]~q ;
wire \F_bht_ptr_nxt[0]~combout ;
wire \M_br_cond_taken_history[1]~q ;
wire \F_bht_ptr_nxt[1]~combout ;
wire \M_br_cond_taken_history[2]~q ;
wire \F_bht_ptr_nxt[2]~combout ;
wire \M_br_cond_taken_history[3]~q ;
wire \F_bht_ptr_nxt[3]~combout ;
wire \M_br_cond_taken_history[4]~q ;
wire \F_bht_ptr_nxt[4]~combout ;
wire \M_br_cond_taken_history[5]~q ;
wire \F_bht_ptr_nxt[5]~combout ;
wire \M_br_cond_taken_history[6]~q ;
wire \F_bht_ptr_nxt[6]~combout ;
wire \M_br_cond_taken_history[7]~q ;
wire \F_bht_ptr_nxt[7]~combout ;
wire \ic_tag_clr_valid_bits_nxt~combout ;
wire \ic_tag_wraddress_nxt~6_combout ;
wire \ic_tag_wraddress_nxt[1]~7_combout ;
wire \ic_tag_wraddress_nxt[2]~8_combout ;
wire \ic_tag_wraddress_nxt[3]~9_combout ;
wire \ic_tag_wraddress_nxt[4]~10_combout ;
wire \ic_tag_wraddress_nxt[5]~11_combout ;
wire \the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[6]~q ;
wire \the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[22]~q ;
wire \the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[7]~q ;
wire \the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[23]~q ;
wire \the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[8]~q ;
wire \the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[24]~q ;
wire \the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[9]~q ;
wire \the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[25]~q ;
wire \the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[15]~q ;
wire \the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[31]~q ;
wire \the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[5]~q ;
wire \the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[21]~q ;
wire \the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[12]~q ;
wire \the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[28]~q ;
wire \the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[11]~q ;
wire \the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[27]~q ;
wire \the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[10]~q ;
wire \the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[26]~q ;
wire \the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[4]~q ;
wire \the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[20]~q ;
wire \the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[3]~q ;
wire \the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[19]~q ;
wire \the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[1]~q ;
wire \the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[17]~q ;
wire \the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[14]~q ;
wire \the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[30]~q ;
wire \the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[2]~q ;
wire \the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[18]~q ;
wire \the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[0]~q ;
wire \the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[16]~q ;
wire \the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[13]~q ;
wire \the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[29]~q ;
wire \E_bht_data[0]~q ;
wire \E_br_mispredict~combout ;
wire \E_bht_ptr[0]~q ;
wire \E_bht_ptr[1]~q ;
wire \E_bht_ptr[2]~q ;
wire \E_bht_ptr[3]~q ;
wire \E_bht_ptr[4]~q ;
wire \E_bht_ptr[5]~q ;
wire \E_bht_ptr[6]~q ;
wire \E_bht_ptr[7]~q ;
wire \E_br_result~2_combout ;
wire \M_br_cond_taken_history[0]~0_combout ;
wire \ic_fill_valid_bits_nxt~0_combout ;
wire \ic_fill_valid_bits_en~combout ;
wire \ic_fill_valid_bits_nxt~1_combout ;
wire \ic_fill_valid_bits_nxt~2_combout ;
wire \ic_fill_valid_bits_nxt~3_combout ;
wire \D_bht_data[0]~q ;
wire \D_bht_ptr[0]~q ;
wire \D_bht_ptr[1]~q ;
wire \D_bht_ptr[2]~q ;
wire \D_bht_ptr[3]~q ;
wire \D_bht_ptr[4]~q ;
wire \D_bht_ptr[5]~q ;
wire \D_bht_ptr[6]~q ;
wire \D_bht_ptr[7]~q ;
wire \ic_fill_valid_bits_nxt~4_combout ;
wire \ic_fill_valid_bits_nxt~5_combout ;
wire \ic_fill_valid_bits_nxt~6_combout ;
wire \ic_fill_valid_bits_nxt~7_combout ;
wire \F_bht_ptr[0]~q ;
wire \F_bht_ptr[1]~q ;
wire \F_bht_ptr[2]~q ;
wire \F_bht_ptr[3]~q ;
wire \F_bht_ptr[4]~q ;
wire \F_bht_ptr[5]~q ;
wire \F_bht_ptr[6]~q ;
wire \F_bht_ptr[7]~q ;
wire \ic_tag_clr_valid_bits~0_combout ;
wire \M_br_mispredict~_wirecell_combout ;
wire \M_sel_data_master~q ;
wire \A_valid_from_M~q ;
wire \D_iw[0]~q ;
wire \D_iw[1]~q ;
wire \D_iw[2]~q ;
wire \D_iw[3]~q ;
wire \D_iw[4]~q ;
wire \Equal95~0_combout ;
wire \D_iw[16]~q ;
wire \D_iw[15]~q ;
wire \D_iw[14]~q ;
wire \D_iw[13]~q ;
wire \D_iw[12]~q ;
wire \D_iw[11]~q ;
wire \D_ctrl_shift_rot~2_combout ;
wire \D_ctrl_late_result~3_combout ;
wire \D_ctrl_illegal~4_combout ;
wire \D_ctrl_illegal~2_combout ;
wire \D_ctrl_flush_pipe_always~2_combout ;
wire \Equal149~6_combout ;
wire \D_ctrl_flush_pipe_always~0_combout ;
wire \D_ctrl_flush_pipe_always~1_combout ;
wire \E_ctrl_flush_pipe_always~q ;
wire \M_ctrl_flush_pipe_always~q ;
wire \A_pipe_flush_nxt~0_combout ;
wire \D_ctrl_cmp~4_combout ;
wire \D_ctrl_alu_force_xor~3_combout ;
wire \D_ctrl_alu_subtract~0_combout ;
wire \D_ctrl_alu_subtract~2_combout ;
wire \D_ctrl_alu_subtract~1_combout ;
wire \E_ctrl_alu_subtract~q ;
wire \Equal149~3_combout ;
wire \Equal149~4_combout ;
wire \Equal95~1_combout ;
wire \Equal95~2_combout ;
wire \Equal95~3_combout ;
wire \Equal95~5_combout ;
wire \D_ctrl_alu_signed_comparison~0_combout ;
wire \D_ctrl_alu_signed_comparison~1_combout ;
wire \E_ctrl_alu_signed_comparison~q ;
wire \D_iw[26]~q ;
wire \D_iw[25]~q ;
wire \D_iw[24]~q ;
wire \D_iw[23]~q ;
wire \D_iw[22]~q ;
wire \Equal304~0_combout ;
wire \F_ctrl_b_is_dst~0_combout ;
wire \D_ctrl_b_is_dst~q ;
wire \D_iw[18]~q ;
wire \F_ctrl_implicit_dst_retaddr~0_combout ;
wire \D_ctrl_implicit_dst_retaddr~q ;
wire \F_ctrl_implicit_dst_eretaddr~1_combout ;
wire \F_ctrl_implicit_dst_eretaddr~2_combout ;
wire \F_ctrl_implicit_dst_eretaddr~0_combout ;
wire \D_ctrl_implicit_dst_eretaddr~q ;
wire \D_dst_regnum[1]~0_combout ;
wire \D_iw[21]~q ;
wire \D_dst_regnum[4]~1_combout ;
wire \F_ctrl_ignore_dst~combout ;
wire \D_ctrl_ignore_dst~q ;
wire \D_iw[17]~q ;
wire \D_dst_regnum[0]~2_combout ;
wire \D_iw[19]~q ;
wire \D_dst_regnum[2]~3_combout ;
wire \D_iw[20]~q ;
wire \D_dst_regnum[3]~4_combout ;
wire \Equal302~0_combout ;
wire \D_wr_dst_reg~combout ;
wire \D_regnum_b_cmp_F~0_combout ;
wire \D_regnum_b_cmp_F~combout ;
wire \E_regnum_b_cmp_D~q ;
wire \A_pipe_flush~q ;
wire \Equal149~0_combout ;
wire \E_ctrl_trap_inst_nxt~combout ;
wire \E_ctrl_trap_inst~q ;
wire \M_exc_trap_inst_pri15~q ;
wire \D_ctrl_unimp_trap~0_combout ;
wire \D_ctrl_unimp_trap~1_combout ;
wire \E_ctrl_unimp_trap~q ;
wire \M_exc_unimp_inst_pri15~q ;
wire \E_iw[15]~q ;
wire \E_iw[14]~q ;
wire \E_iw[12]~q ;
wire \E_iw[11]~q ;
wire \E_iw[16]~q ;
wire \E_iw[13]~q ;
wire \E_iw[1]~q ;
wire \E_iw[2]~q ;
wire \E_iw[0]~q ;
wire \E_iw[5]~q ;
wire \E_iw[4]~q ;
wire \E_iw[3]~q ;
wire \Equal239~0_combout ;
wire \E_op_rdctl~0_combout ;
wire \E_op_break~combout ;
wire \M_exc_break_inst_pri15~q ;
wire \D_ctrl_illegal~0_combout ;
wire \D_ctrl_illegal~3_combout ;
wire \D_ctrl_illegal~1_combout ;
wire \E_ctrl_illegal~q ;
wire \M_exc_illegal_inst_pri15~q ;
wire \M_exc_any~0_combout ;
wire \E_wr_dst_reg_from_D~q ;
wire \E_wr_dst_reg~combout ;
wire \M_wr_dst_reg_from_E~q ;
wire \M_wr_dst_reg~0_combout ;
wire \A_wr_dst_reg_from_M~q ;
wire \A_wr_dst_reg~0_combout ;
wire \M_exc_break~0_combout ;
wire \A_exc_break~q ;
wire \E_dst_regnum[0]~q ;
wire \M_dst_regnum[0]~q ;
wire \A_dst_regnum_from_M[0]~q ;
wire \A_dst_regnum~0_combout ;
wire \E_dst_regnum[1]~q ;
wire \M_dst_regnum[1]~q ;
wire \A_dst_regnum_from_M[1]~q ;
wire \A_dst_regnum~1_combout ;
wire \E_dst_regnum[2]~q ;
wire \M_dst_regnum[2]~q ;
wire \A_dst_regnum_from_M[2]~q ;
wire \A_dst_regnum~2_combout ;
wire \A_regnum_b_cmp_F~0_combout ;
wire \E_dst_regnum[3]~q ;
wire \M_dst_regnum[3]~q ;
wire \A_dst_regnum_from_M[3]~q ;
wire \A_dst_regnum~3_combout ;
wire \E_dst_regnum[4]~q ;
wire \M_dst_regnum[4]~q ;
wire \A_dst_regnum_from_M[4]~q ;
wire \A_dst_regnum~4_combout ;
wire \A_regnum_b_cmp_F~1_combout ;
wire \A_regnum_b_cmp_F~combout ;
wire \M_regnum_b_cmp_F~0_combout ;
wire \M_regnum_b_cmp_F~1_combout ;
wire \M_regnum_b_cmp_F~combout ;
wire \E_regnum_b_cmp_F~0_combout ;
wire \E_regnum_b_cmp_F~1_combout ;
wire \E_regnum_b_cmp_F~combout ;
wire \M_regnum_b_cmp_D~q ;
wire \A_regnum_b_cmp_D~q ;
wire \W_regnum_b_cmp_D~q ;
wire \D_src2_reg[0]~0_combout ;
wire \D_src2_reg[0]~4_combout ;
wire \D_src2_reg[0]~1_combout ;
wire \D_src2_reg[0]~5_combout ;
wire \D_src2_reg[0]~6_combout ;
wire \F_ctrl_src2_choose_imm~1_combout ;
wire \F_ctrl_src2_choose_imm~0_combout ;
wire \D_ctrl_src2_choose_imm~q ;
wire \D_ctrl_logic~0_combout ;
wire \D_ctrl_logic~1_combout ;
wire \E_ctrl_logic~q ;
wire \Equal95~4_combout ;
wire \D_ctrl_retaddr~1_combout ;
wire \D_ctrl_retaddr~0_combout ;
wire \E_ctrl_retaddr~q ;
wire \E_alu_result~0_combout ;
wire \D_src2_reg[0]~2_combout ;
wire \D_logic_op_raw[1]~1_combout ;
wire \D_ctrl_alu_force_xor~1_combout ;
wire \Equal149~5_combout ;
wire \Equal149~1_combout ;
wire \Equal149~2_combout ;
wire \D_ctrl_alu_force_xor~0_combout ;
wire \D_ctrl_alu_force_xor~2_combout ;
wire \D_logic_op[1]~0_combout ;
wire \E_logic_op[1]~q ;
wire \D_logic_op_raw[0]~0_combout ;
wire \D_logic_op[0]~1_combout ;
wire \E_logic_op[0]~q ;
wire \E_alu_result~10_combout ;
wire \E_alu_result[31]~combout ;
wire \M_alu_result[31]~q ;
wire \Equal219~0_combout ;
wire \Equal219~1_combout ;
wire \M_ctrl_ld32~q ;
wire \A_ctrl_ld32~q ;
wire \d_readdata_d1[31]~q ;
wire \M_alu_result[1]~q ;
wire \d_readdata_d1[1]~q ;
wire \d_readdata_d1[17]~q ;
wire \d_readdata_d1[9]~q ;
wire \d_readdata_d1[25]~q ;
wire \Equal212~0_combout ;
wire \Equal212~1_combout ;
wire \M_ctrl_ld8~q ;
wire \Equal215~0_combout ;
wire \M_ctrl_ld16~q ;
wire \M_ld_align_sh16~0_combout ;
wire \A_ld_align_sh16~q ;
wire \F_ctrl_hi_imm16~0_combout ;
wire \D_ctrl_hi_imm16~q ;
wire \D_ctrl_shift_right_arith~0_combout ;
wire \E_src2[1]~0_combout ;
wire \D_iw[6]~q ;
wire \d_readdata_d1[0]~q ;
wire \d_readdata_d1[16]~q ;
wire \d_readdata_d1[8]~q ;
wire \d_readdata_d1[24]~q ;
wire \A_slow_inst_result_nxt[0]~0_combout ;
wire \D_ctrl_ld~0_combout ;
wire \E_ctrl_ld~q ;
wire \M_ctrl_ld~q ;
wire \A_ctrl_ld~q ;
wire \A_slow_inst_result[0]~q ;
wire \D_ctrl_shift_right_arith~1_combout ;
wire \D_ctrl_shift_right_arith~2_combout ;
wire \E_ctrl_shift_right_arith~q ;
wire \E_rot_fill_bit~0_combout ;
wire \M_rot_fill_bit~q ;
wire \M_alu_result[3]~q ;
wire \d_readdata_d1[3]~q ;
wire \d_readdata_d1[19]~q ;
wire \d_readdata_d1[11]~q ;
wire \d_readdata_d1[27]~q ;
wire \A_slow_inst_result_nxt[3]~3_combout ;
wire \A_slow_inst_result[3]~q ;
wire \M_alu_result[4]~q ;
wire \d_readdata_d1[4]~q ;
wire \d_readdata_d1[20]~q ;
wire \d_readdata_d1[12]~q ;
wire \d_readdata_d1[28]~q ;
wire \A_slow_inst_result_nxt[4]~4_combout ;
wire \A_slow_inst_result[4]~q ;
wire \M_alu_result[2]~q ;
wire \d_readdata_d1[2]~q ;
wire \d_readdata_d1[18]~q ;
wire \d_readdata_d1[10]~q ;
wire \d_readdata_d1[26]~q ;
wire \A_slow_inst_result_nxt[2]~2_combout ;
wire \A_slow_inst_result[2]~q ;
wire \E_ctrl_shift_rot_right~q ;
wire \E_rot_mask[2]~2_combout ;
wire \M_rot_mask[2]~q ;
wire \D_src2_reg[0]~7_combout ;
wire \D_src2_reg[0]~8_combout ;
wire \M_ctrl_ld8_ld16~q ;
wire \M_ld_align_byte2_byte3_fill~combout ;
wire \A_ld_align_byte2_byte3_fill~q ;
wire \d_readdata_d1[22]~q ;
wire \A_slow_inst_result_nxt[22]~35_combout ;
wire \A_slow_inst_result_nxt[22]~8_combout ;
wire \A_slow_inst_result[22]~q ;
wire \E_rot_mask[6]~6_combout ;
wire \M_rot_mask[6]~q ;
wire \D_ctrl_rot~0_combout ;
wire \E_ctrl_rot~q ;
wire \D_ctrl_shift_rot_left~0_combout ;
wire \E_ctrl_shift_rot_left~q ;
wire \E_rot_pass2~0_combout ;
wire \M_rot_pass2~q ;
wire \E_rot_sel_fill2~0_combout ;
wire \M_rot_sel_fill2~q ;
wire \A_slow_inst_result_nxt[18]~32_combout ;
wire \A_slow_inst_result_nxt[18]~21_combout ;
wire \A_slow_inst_result[18]~q ;
wire \M_ld_align_byte1_fill~0_combout ;
wire \A_ld_align_byte1_fill~q ;
wire \A_slow_inst_result[9]~1_combout ;
wire \d_readdata_d1[14]~q ;
wire \d_readdata_d1[30]~q ;
wire \A_slow_inst_result[9]~0_combout ;
wire \A_slow_inst_result_nxt[14]~46_combout ;
wire \A_slow_inst_result_nxt[14]~48_combout ;
wire \A_slow_inst_result[14]~q ;
wire \E_rot_pass1~0_combout ;
wire \M_rot_pass1~q ;
wire \E_rot_sel_fill1~0_combout ;
wire \M_rot_sel_fill1~q ;
wire \A_slow_inst_result_nxt[10]~42_combout ;
wire \A_slow_inst_result_nxt[10]~72_combout ;
wire \A_slow_inst_result[10]~q ;
wire \d_readdata_d1[6]~q ;
wire \A_slow_inst_result_nxt[6]~6_combout ;
wire \A_slow_inst_result[6]~q ;
wire \E_compare_op[0]~q ;
wire \E_logic_result[3]~0_combout ;
wire \Equal316~0_combout ;
wire \Equal316~1_combout ;
wire \Equal316~2_combout ;
wire \d_readdata_d1[7]~q ;
wire \d_readdata_d1[23]~q ;
wire \d_readdata_d1[15]~q ;
wire \A_slow_inst_result_nxt[7]~7_combout ;
wire \A_slow_inst_result[7]~q ;
wire \E_rot_mask[7]~7_combout ;
wire \M_rot_mask[7]~q ;
wire \Add10~0_combout ;
wire \E_rot_step1[3]~25_combout ;
wire \d_readdata_d1[5]~q ;
wire \d_readdata_d1[21]~q ;
wire \d_readdata_d1[13]~q ;
wire \d_readdata_d1[29]~q ;
wire \A_slow_inst_result_nxt[5]~5_combout ;
wire \A_slow_inst_result[5]~q ;
wire \E_rot_mask[5]~5_combout ;
wire \M_rot_mask[5]~q ;
wire \E_rot_step1[1]~9_combout ;
wire \Add9~134_cout ;
wire \Add9~66 ;
wire \Add9~70 ;
wire \Add9~58 ;
wire \Add9~54 ;
wire \Add9~2 ;
wire \Add9~5_sumout ;
wire \E_alu_result~4_combout ;
wire \D_pc[3]~q ;
wire \D_iw[9]~q ;
wire \Equal95~6_combout ;
wire \F_ctrl_br~0_combout ;
wire \D_ctrl_br~q ;
wire \D_bht_data[1]~q ;
wire \F_ctrl_br_uncond~0_combout ;
wire \D_ctrl_br_uncond~q ;
wire \D_br_pred_taken~0_combout ;
wire \F_older_non_sequential~0_combout ;
wire \E_ctrl_jmp_indirect_nxt~0_combout ;
wire \E_valid_jmp_indirect~0_combout ;
wire \E_valid_jmp_indirect~q ;
wire \D_pc[2]~q ;
wire \D_pc[1]~q ;
wire \D_pc[0]~q ;
wire \Add3~1_sumout ;
wire \Add0~1_sumout ;
wire \D_br_taken_waddr_partial[0]~q ;
wire \D_kill~q ;
wire \F_ic_tag_rd_addr_nxt[3]~1_combout ;
wire \F_ic_data_rd_addr_nxt[0]~0_combout ;
wire \E_pc[0]~q ;
wire \M_pc_plus_one[0]~0_combout ;
wire \M_pc_plus_one[0]~q ;
wire \M_target_pcb[2]~q ;
wire \E_ctrl_jmp_indirect~q ;
wire \M_ctrl_jmp_indirect~q ;
wire \A_pipe_flush_waddr_nxt~0_combout ;
wire \A_pipe_flush_waddr[0]~q ;
wire \D_pc_plus_one[0]~q ;
wire \E_ctrl_br_cond_nxt~0_combout ;
wire \D_br_pred_not_taken~combout ;
wire \E_extra_pc[0]~q ;
wire \M_pipe_flush_waddr[0]~q ;
wire \F_ic_tag_rd_addr_nxt[3]~2_combout ;
wire \F_ic_tag_rd_addr_nxt[3]~3_combout ;
wire \F_ic_data_rd_addr_nxt[0]~1_combout ;
wire \F_pc[0]~q ;
wire \Add3~2 ;
wire \Add3~5_sumout ;
wire \Add0~2 ;
wire \Add0~5_sumout ;
wire \D_br_taken_waddr_partial[1]~q ;
wire \D_iw[7]~q ;
wire \F_ic_data_rd_addr_nxt[1]~2_combout ;
wire \E_pc[1]~q ;
wire \Add7~1_sumout ;
wire \M_pc_plus_one[1]~q ;
wire \M_target_pcb[3]~q ;
wire \A_pipe_flush_waddr_nxt~1_combout ;
wire \A_pipe_flush_waddr[1]~q ;
wire \D_pc_plus_one[1]~q ;
wire \E_extra_pc[1]~q ;
wire \M_pipe_flush_waddr[1]~q ;
wire \F_ic_data_rd_addr_nxt[1]~3_combout ;
wire \F_pc[1]~q ;
wire \Add3~6 ;
wire \Add3~9_sumout ;
wire \Add0~6 ;
wire \Add0~9_sumout ;
wire \D_br_taken_waddr_partial[2]~q ;
wire \D_iw[8]~q ;
wire \F_ic_data_rd_addr_nxt[2]~4_combout ;
wire \E_pc[2]~q ;
wire \Add7~2 ;
wire \Add7~5_sumout ;
wire \M_pc_plus_one[2]~q ;
wire \M_target_pcb[4]~q ;
wire \A_pipe_flush_waddr_nxt~2_combout ;
wire \A_pipe_flush_waddr[2]~q ;
wire \D_pc_plus_one[2]~q ;
wire \E_extra_pc[2]~q ;
wire \M_pipe_flush_waddr[2]~q ;
wire \F_ic_data_rd_addr_nxt[2]~5_combout ;
wire \F_pc[2]~q ;
wire \F_ic_valid~4_combout ;
wire \F_ic_valid~0_combout ;
wire \D_pc[14]~q ;
wire \D_pc[13]~q ;
wire \D_pc[12]~q ;
wire \D_pc[11]~q ;
wire \D_pc[10]~q ;
wire \D_pc[9]~q ;
wire \D_pc[8]~q ;
wire \D_pc[7]~q ;
wire \D_pc[6]~q ;
wire \D_pc[5]~q ;
wire \D_pc[4]~q ;
wire \Add3~10 ;
wire \Add3~14 ;
wire \Add3~17_sumout ;
wire \Add0~10 ;
wire \Add0~14 ;
wire \Add0~17_sumout ;
wire \D_br_taken_waddr_partial[4]~q ;
wire \D_iw[10]~q ;
wire \F_ic_tag_rd_addr_nxt[1]~6_combout ;
wire \E_pc[4]~q ;
wire \E_pc[3]~q ;
wire \Add7~6 ;
wire \Add7~10 ;
wire \Add7~13_sumout ;
wire \M_pc_plus_one[4]~q ;
wire \M_target_pcb[6]~q ;
wire \A_pipe_flush_waddr_nxt~4_combout ;
wire \A_pipe_flush_waddr[4]~q ;
wire \D_pc_plus_one[4]~q ;
wire \E_extra_pc[4]~q ;
wire \M_pipe_flush_waddr[4]~q ;
wire \F_ic_tag_rd_addr_nxt[1]~7_combout ;
wire \F_pc[4]~q ;
wire \Add3~18 ;
wire \Add3~21_sumout ;
wire \Add0~18 ;
wire \Add0~21_sumout ;
wire \D_br_taken_waddr_partial[5]~q ;
wire \F_ic_tag_rd_addr_nxt[2]~8_combout ;
wire \E_pc[5]~q ;
wire \Add7~14 ;
wire \Add7~17_sumout ;
wire \M_pc_plus_one[5]~q ;
wire \M_target_pcb[7]~q ;
wire \A_pipe_flush_waddr_nxt~5_combout ;
wire \A_pipe_flush_waddr[5]~q ;
wire \D_pc_plus_one[5]~q ;
wire \E_extra_pc[5]~q ;
wire \M_pipe_flush_waddr[5]~q ;
wire \F_ic_tag_rd_addr_nxt[2]~9_combout ;
wire \F_pc[5]~q ;
wire \Add3~22 ;
wire \Add3~25_sumout ;
wire \Add0~22 ;
wire \Add0~33_sumout ;
wire \D_br_taken_waddr_partial[6]~q ;
wire \F_ic_tag_rd_addr_nxt[3]~10_combout ;
wire \A_slow_inst_result_nxt[8]~40_combout ;
wire \A_slow_inst_result_nxt[8]~68_combout ;
wire \A_slow_inst_result[8]~q ;
wire \E_rot_mask[0]~0_combout ;
wire \M_rot_mask[0]~q ;
wire \E_rot_step1[4]~6_combout ;
wire \E_rot_step1[8]~7_combout ;
wire \Add10~1_combout ;
wire \M_rot_prestep2[8]~q ;
wire \E_rot_step1[28]~0_combout ;
wire \E_rot_step1[0]~1_combout ;
wire \M_rot_prestep2[0]~q ;
wire \A_slow_inst_result_nxt[20]~34_combout ;
wire \A_slow_inst_result_nxt[20]~17_combout ;
wire \A_slow_inst_result[20]~q ;
wire \A_slow_inst_result_nxt[16]~29_combout ;
wire \A_slow_inst_result_nxt[16]~22_combout ;
wire \A_slow_inst_result[16]~q ;
wire \A_slow_inst_result_nxt[12]~44_combout ;
wire \A_slow_inst_result_nxt[12]~56_combout ;
wire \A_slow_inst_result[12]~q ;
wire \M_rot_prestep2[12]~q ;
wire \M_rot_prestep2[4]~q ;
wire \A_slow_inst_result_nxt[21]~27_combout ;
wire \A_slow_inst_result_nxt[21]~13_combout ;
wire \A_slow_inst_result[21]~q ;
wire \A_slow_inst_result_nxt[17]~30_combout ;
wire \A_slow_inst_result_nxt[17]~19_combout ;
wire \A_slow_inst_result[17]~q ;
wire \E_rot_mask[1]~1_combout ;
wire \M_rot_mask[1]~q ;
wire \A_slow_inst_result_nxt[13]~45_combout ;
wire \A_slow_inst_result_nxt[13]~52_combout ;
wire \A_slow_inst_result[13]~q ;
wire \A_slow_inst_result_nxt[9]~41_combout ;
wire \A_slow_inst_result_nxt[9]~64_combout ;
wire \A_slow_inst_result[9]~q ;
wire \M_rot_prestep2[9]~q ;
wire \E_rot_step1[29]~8_combout ;
wire \M_rot_prestep2[1]~q ;
wire \A_slow_inst_result_nxt[19]~33_combout ;
wire \A_slow_inst_result_nxt[19]~18_combout ;
wire \A_slow_inst_result[19]~q ;
wire \E_rot_mask[3]~3_combout ;
wire \M_rot_mask[3]~q ;
wire \A_slow_inst_result_nxt[15]~47_combout ;
wire \A_slow_inst_result_nxt[15]~60_combout ;
wire \A_slow_inst_result[15]~q ;
wire \A_slow_inst_result_nxt[11]~43_combout ;
wire \A_slow_inst_result_nxt[11]~76_combout ;
wire \A_slow_inst_result[11]~q ;
wire \M_rot_prestep2[11]~q ;
wire \E_rot_step1[31]~24_combout ;
wire \M_rot_prestep2[3]~q ;
wire \E_rot_step1[23]~26_combout ;
wire \E_rot_step1[27]~27_combout ;
wire \M_rot_prestep2[27]~q ;
wire \Add10~2_combout ;
wire \M_rot_rn[3]~q ;
wire \Add10~3_combout ;
wire \M_rot_rn[4]~q ;
wire \M_rot[3]~14_combout ;
wire \A_shift_rot_result~14_combout ;
wire \A_shift_rot_result[11]~q ;
wire \E_pc[9]~q ;
wire \E_pc[8]~q ;
wire \E_pc[7]~q ;
wire \E_pc[6]~q ;
wire \Add7~18 ;
wire \Add7~30 ;
wire \Add7~34 ;
wire \Add7~26 ;
wire \Add7~21_sumout ;
wire \M_pc_plus_one[9]~q ;
wire \E_op_rdctl~1_combout ;
wire \E_op_rdctl~combout ;
wire \M_ctrl_rd_ctl_reg~q ;
wire \A_inst_result[9]~0_combout ;
wire \A_inst_result[11]~q ;
wire \A_mul_cell_p1[11]~q ;
wire \Equal95~7_combout ;
wire \D_ctrl_late_result~2_combout ;
wire \D_ctrl_mul_lsw~0_combout ;
wire \E_ctrl_mul_lsw~q ;
wire \M_ctrl_mul_lsw~q ;
wire \A_ctrl_mul_lsw~q ;
wire \D_ctrl_shift_rot~0_combout ;
wire \E_ctrl_shift_rot~q ;
wire \M_ctrl_shift_rot~q ;
wire \A_ctrl_shift_rot~q ;
wire \A_wr_data_unfiltered[15]~0_combout ;
wire \A_slow_inst_sel_nxt~0_combout ;
wire \A_slow_inst_sel~q ;
wire \A_wr_data_unfiltered[15]~1_combout ;
wire \A_wr_data_unfiltered[11]~16_combout ;
wire \W_wr_data[11]~q ;
wire \D_src2_reg[11]~38_combout ;
wire \D_src2_reg[11]~39_combout ;
wire \E_src2[5]~2_combout ;
wire \E_src2[11]~q ;
wire \Add9~46 ;
wire \Add9~10 ;
wire \Add9~42 ;
wire \Add9~38 ;
wire \Add9~33_sumout ;
wire \E_alu_result~11_combout ;
wire \D_pc_plus_one[9]~q ;
wire \E_extra_pc[9]~q ;
wire \E_alu_result[11]~combout ;
wire \M_alu_result[11]~q ;
wire \F_ctrl_a_not_src~0_combout ;
wire \D_ctrl_a_not_src~q ;
wire \E_regnum_a_cmp_F~0_combout ;
wire \E_regnum_a_cmp_F~1_combout ;
wire \E_regnum_a_cmp_F~combout ;
wire \D_regnum_a_cmp_F~0_combout ;
wire \D_regnum_a_cmp_F~combout ;
wire \E_regnum_a_cmp_D~q ;
wire \M_regnum_a_cmp_D~q ;
wire \A_regnum_a_cmp_F~0_combout ;
wire \A_regnum_a_cmp_F~1_combout ;
wire \A_regnum_a_cmp_F~combout ;
wire \M_regnum_a_cmp_F~0_combout ;
wire \M_regnum_a_cmp_F~1_combout ;
wire \M_regnum_a_cmp_F~combout ;
wire \A_regnum_a_cmp_D~q ;
wire \W_regnum_a_cmp_D~q ;
wire \E_src1[26]~0_combout ;
wire \E_src1[26]~1_combout ;
wire \D_src1_reg[11]~10_combout ;
wire \D_iw[31]~q ;
wire \D_iw[30]~q ;
wire \D_iw[29]~q ;
wire \D_iw[28]~q ;
wire \D_iw[27]~q ;
wire \Equal303~0_combout ;
wire \D_src1_hazard_E~combout ;
wire \E_src1[11]~q ;
wire \E_rot_step1[11]~31_combout ;
wire \M_rot_prestep2[15]~q ;
wire \M_rot_prestep2[31]~q ;
wire \E_rot_step1[19]~29_combout ;
wire \M_rot_prestep2[23]~q ;
wire \M_rot[7]~27_combout ;
wire \A_shift_rot_result~27_combout ;
wire \A_shift_rot_result[15]~q ;
wire \E_pc[13]~q ;
wire \E_pc[12]~q ;
wire \E_pc[11]~q ;
wire \E_pc[10]~q ;
wire \Add7~22 ;
wire \Add7~46 ;
wire \Add7~50 ;
wire \Add7~54 ;
wire \Add7~41_sumout ;
wire \M_pc_plus_one[13]~q ;
wire \A_inst_result[15]~q ;
wire \A_mul_cell_p1[15]~q ;
wire \A_wr_data_unfiltered[15]~29_combout ;
wire \W_wr_data[15]~q ;
wire \D_src2_reg[15]~62_combout ;
wire \D_src2_reg[15]~63_combout ;
wire \E_src2[15]~q ;
wire \Add9~34 ;
wire \Add9~30 ;
wire \Add9~26 ;
wire \Add9~22 ;
wire \Add9~17_sumout ;
wire \E_alu_result~20_combout ;
wire \E_extra_pc[13]~q ;
wire \E_alu_result[15]~combout ;
wire \M_alu_result[15]~q ;
wire \D_src1_reg[15]~27_combout ;
wire \E_src1[15]~q ;
wire \E_rot_step1[15]~28_combout ;
wire \M_rot_prestep2[19]~q ;
wire \M_rot[3]~22_combout ;
wire \A_shift_rot_result~22_combout ;
wire \A_shift_rot_result[19]~q ;
wire \A_inst_result[26]~1_combout ;
wire \A_inst_result[19]~q ;
wire \Add11~58 ;
wire \Add11~46 ;
wire \Add11~54 ;
wire \Add11~41_sumout ;
wire \A_mul_s1[3]~q ;
wire \A_mul_cell_p3[3]~q ;
wire \Add11~53_sumout ;
wire \A_mul_s1[2]~q ;
wire \A_mul_cell_p3[2]~q ;
wire \Add11~45_sumout ;
wire \A_mul_s1[1]~q ;
wire \A_mul_cell_p3[1]~q ;
wire \Add11~57_sumout ;
wire \A_mul_s1[0]~q ;
wire \A_mul_cell_p3[0]~q ;
wire \Add12~58 ;
wire \Add12~46 ;
wire \Add12~54 ;
wire \Add12~41_sumout ;
wire \A_wr_data_unfiltered[19]~24_combout ;
wire \W_wr_data[19]~q ;
wire \D_src2_reg[19]~55_combout ;
wire \Add9~18 ;
wire \Add9~14 ;
wire \Add9~118 ;
wire \Add9~126 ;
wire \Add9~113_sumout ;
wire \Equal0~0_combout ;
wire \F_ctrl_unsigned_lo_imm16~1_combout ;
wire \F_ctrl_unsigned_lo_imm16~0_combout ;
wire \D_ctrl_unsigned_lo_imm16~q ;
wire \D_src2[19]~37_combout ;
wire \D_src2[19]~38_combout ;
wire \D_src2[19]~20_combout ;
wire \E_src2[30]~1_combout ;
wire \E_src2[19]~q ;
wire \E_logic_result[19]~10_combout ;
wire \E_alu_result[19]~combout ;
wire \M_alu_result[19]~q ;
wire \D_src1_reg[19]~21_combout ;
wire \E_src1[19]~q ;
wire \E_rot_step1[21]~10_combout ;
wire \E_rot_step1[25]~11_combout ;
wire \M_rot_prestep2[25]~q ;
wire \M_rot[1]~19_combout ;
wire \A_shift_rot_result~19_combout ;
wire \A_shift_rot_result[9]~q ;
wire \Add7~33_sumout ;
wire \M_pc_plus_one[7]~q ;
wire \A_inst_result[9]~q ;
wire \A_mul_cell_p1[9]~q ;
wire \A_wr_data_unfiltered[9]~21_combout ;
wire \W_wr_data[9]~q ;
wire \D_src2_reg[9]~50_combout ;
wire \D_src2_reg[9]~51_combout ;
wire \E_src2[9]~q ;
wire \Add9~41_sumout ;
wire \E_alu_result~16_combout ;
wire \D_pc_plus_one[7]~q ;
wire \E_extra_pc[7]~q ;
wire \E_alu_result[9]~combout ;
wire \M_alu_result[9]~q ;
wire \D_src1_reg[9]~15_combout ;
wire \E_src1[9]~q ;
wire \E_rot_step1[9]~15_combout ;
wire \M_rot_prestep2[13]~q ;
wire \M_rot_prestep2[29]~q ;
wire \M_rot[5]~29_combout ;
wire \A_shift_rot_result~29_combout ;
wire \A_shift_rot_result[13]~q ;
wire \Add7~49_sumout ;
wire \M_pc_plus_one[11]~q ;
wire \A_inst_result[13]~q ;
wire \A_mul_cell_p1[13]~q ;
wire \A_wr_data_unfiltered[13]~31_combout ;
wire \W_wr_data[13]~q ;
wire \D_src2_reg[13]~66_combout ;
wire \D_src2_reg[13]~67_combout ;
wire \E_src2[13]~q ;
wire \Add9~25_sumout ;
wire \E_alu_result~22_combout ;
wire \E_extra_pc[11]~q ;
wire \E_alu_result[13]~combout ;
wire \M_alu_result[13]~q ;
wire \D_src1_reg[13]~29_combout ;
wire \E_src1[13]~q ;
wire \E_rot_step1[13]~12_combout ;
wire \M_rot_prestep2[17]~q ;
wire \M_rot[1]~23_combout ;
wire \A_shift_rot_result~23_combout ;
wire \A_shift_rot_result[17]~q ;
wire \A_inst_result[17]~q ;
wire \Add12~45_sumout ;
wire \A_wr_data_unfiltered[17]~25_combout ;
wire \W_wr_data[17]~q ;
wire \D_src2_reg[17]~56_combout ;
wire \Add9~117_sumout ;
wire \D_src2[17]~33_combout ;
wire \D_src2[17]~34_combout ;
wire \D_src2[17]~21_combout ;
wire \E_src2[17]~q ;
wire \E_logic_result[17]~4_combout ;
wire \E_alu_result[17]~combout ;
wire \M_alu_result[17]~q ;
wire \D_src1_reg[17]~22_combout ;
wire \E_src1[17]~q ;
wire \E_rot_step1[17]~13_combout ;
wire \M_rot_prestep2[21]~q ;
wire \M_rot[5]~13_combout ;
wire \A_shift_rot_result~13_combout ;
wire \A_shift_rot_result[21]~q ;
wire \A_inst_result[21]~q ;
wire \Add11~42 ;
wire \Add11~38 ;
wire \Add11~21_sumout ;
wire \A_mul_s1[5]~q ;
wire \A_mul_cell_p3[5]~q ;
wire \Add11~37_sumout ;
wire \A_mul_s1[4]~q ;
wire \A_mul_cell_p3[4]~q ;
wire \Add12~42 ;
wire \Add12~38 ;
wire \Add12~21_sumout ;
wire \A_wr_data_unfiltered[21]~15_combout ;
wire \W_wr_data[21]~q ;
wire \D_src2_reg[21]~37_combout ;
wire \Add9~114 ;
wire \Add9~110 ;
wire \Add9~93_sumout ;
wire \D_src2[21]~29_combout ;
wire \D_src2[21]~30_combout ;
wire \D_src2[21]~11_combout ;
wire \E_src2[21]~q ;
wire \E_logic_result[21]~8_combout ;
wire \E_alu_result[21]~combout ;
wire \M_alu_result[21]~q ;
wire \D_src1_reg[21]~9_combout ;
wire \E_src1[21]~q ;
wire \E_rot_step1[24]~3_combout ;
wire \M_rot_prestep2[28]~q ;
wire \M_rot[4]~28_combout ;
wire \A_shift_rot_result~28_combout ;
wire \A_shift_rot_result[12]~q ;
wire \Add7~45_sumout ;
wire \M_pc_plus_one[10]~q ;
wire \A_inst_result[12]~q ;
wire \A_mul_cell_p1[12]~q ;
wire \A_wr_data_unfiltered[12]~30_combout ;
wire \W_wr_data[12]~q ;
wire \D_src2_reg[12]~64_combout ;
wire \D_src2_reg[12]~65_combout ;
wire \E_src2[12]~q ;
wire \Add9~29_sumout ;
wire \E_alu_result~21_combout ;
wire \E_extra_pc[10]~q ;
wire \E_alu_result[12]~combout ;
wire \M_alu_result[12]~q ;
wire \D_src1_reg[12]~28_combout ;
wire \E_src1[12]~q ;
wire \E_rot_step1[12]~4_combout ;
wire \M_rot_prestep2[16]~q ;
wire \M_rot[0]~26_combout ;
wire \A_shift_rot_result~26_combout ;
wire \A_shift_rot_result[16]~q ;
wire \E_pc[14]~q ;
wire \Add7~42 ;
wire \Add7~37_sumout ;
wire \M_pc_plus_one[14]~q ;
wire \E_iw[9]~q ;
wire \E_iw[7]~q ;
wire \E_iw[6]~q ;
wire \E_iw[10]~q ;
wire \E_iw[8]~q ;
wire \M_control_reg_rddata[16]~0_combout ;
wire \M_iw[7]~q ;
wire \A_iw[7]~q ;
wire \M_iw[6]~q ;
wire \A_iw[6]~q ;
wire \M_iw[10]~q ;
wire \A_iw[10]~q ;
wire \M_iw[9]~q ;
wire \A_iw[9]~q ;
wire \M_iw[8]~q ;
wire \A_iw[8]~q ;
wire \E_op_wrctl~combout ;
wire \M_ctrl_wrctl_inst~q ;
wire \A_ctrl_wrctl_inst~q ;
wire \A_wrctl_status~0_combout ;
wire \W_ienable_reg_irq1_nxt~0_combout ;
wire \W_ienable_reg_irq16~q ;
wire \W_ipending_reg_irq16_nxt~0_combout ;
wire \W_ipending_reg_irq16~q ;
wire \Equal324~0_combout ;
wire \E_control_reg_rddata[1]~0_combout ;
wire \D_control_reg_rddata_muxed[16]~3_combout ;
wire \E_control_reg_rddata[16]~q ;
wire \E_control_reg_rddata_muxed[16]~5_combout ;
wire \M_control_reg_rddata[16]~q ;
wire \M_inst_result[16]~5_combout ;
wire \A_inst_result[16]~q ;
wire \Add12~57_sumout ;
wire \A_wr_data_unfiltered[16]~28_combout ;
wire \W_wr_data[16]~q ;
wire \D_src2_reg[16]~61_combout ;
wire \E_logic_result[16]~12_combout ;
wire \E_extra_pc[14]~q ;
wire \E_alu_result[16]~19_combout ;
wire \D_src2[16]~31_combout ;
wire \D_src2[16]~32_combout ;
wire \D_src2[16]~26_combout ;
wire \E_src2[16]~q ;
wire \Add9~13_sumout ;
wire \E_alu_result[16]~combout ;
wire \M_alu_result[16]~q ;
wire \D_src1_reg[16]~26_combout ;
wire \E_src1[16]~q ;
wire \E_rot_step1[16]~5_combout ;
wire \M_rot_prestep2[20]~q ;
wire \M_rot[4]~21_combout ;
wire \A_shift_rot_result~21_combout ;
wire \A_shift_rot_result[20]~q ;
wire \A_inst_result[20]~q ;
wire \Add12~37_sumout ;
wire \A_wr_data_unfiltered[20]~23_combout ;
wire \W_wr_data[20]~q ;
wire \D_src2_reg[20]~54_combout ;
wire \Add9~109_sumout ;
wire \D_src2[20]~39_combout ;
wire \D_src2[20]~40_combout ;
wire \D_src2[20]~19_combout ;
wire \E_src2[20]~q ;
wire \E_logic_result[20]~9_combout ;
wire \E_alu_result[20]~combout ;
wire \M_alu_result[20]~q ;
wire \D_src1_reg[20]~20_combout ;
wire \E_src1[20]~q ;
wire \E_rot_step1[20]~2_combout ;
wire \M_rot_prestep2[24]~q ;
wire \M_rot[0]~18_combout ;
wire \A_shift_rot_result~18_combout ;
wire \A_shift_rot_result[8]~q ;
wire \Add7~29_sumout ;
wire \M_pc_plus_one[6]~q ;
wire \A_inst_result[8]~q ;
wire \A_mul_cell_p1[8]~q ;
wire \A_wr_data_unfiltered[8]~20_combout ;
wire \W_wr_data[8]~q ;
wire \D_src2_reg[8]~48_combout ;
wire \D_src2_reg[8]~49_combout ;
wire \E_src2[8]~q ;
wire \Add9~9_sumout ;
wire \E_alu_result~15_combout ;
wire \D_pc_plus_one[6]~q ;
wire \E_extra_pc[6]~q ;
wire \E_alu_result[8]~combout ;
wire \M_alu_result[8]~q ;
wire \D_src1_reg[8]~14_combout ;
wire \E_src1[8]~q ;
wire \M_target_pcb[8]~q ;
wire \A_pipe_flush_waddr_nxt~6_combout ;
wire \A_pipe_flush_waddr[6]~q ;
wire \M_pipe_flush_waddr[6]~q ;
wire \F_ic_tag_rd_addr_nxt[3]~11_combout ;
wire \F_pc[6]~q ;
wire \Add3~26 ;
wire \Add3~29_sumout ;
wire \Add0~34 ;
wire \Add0~37_sumout ;
wire \D_br_taken_waddr_partial[7]~q ;
wire \F_ic_tag_rd_addr_nxt[4]~12_combout ;
wire \M_target_pcb[9]~q ;
wire \A_pipe_flush_waddr_nxt~7_combout ;
wire \A_pipe_flush_waddr[7]~q ;
wire \M_pipe_flush_waddr[7]~q ;
wire \F_ic_tag_rd_addr_nxt[4]~13_combout ;
wire \F_pc[7]~q ;
wire \Add3~30 ;
wire \Add3~33_sumout ;
wire \Add0~38 ;
wire \Add0~29_sumout ;
wire \D_br_taken_waddr_partial[8]~q ;
wire \F_ic_tag_rd_addr_nxt[5]~14_combout ;
wire \Add7~25_sumout ;
wire \M_pc_plus_one[8]~q ;
wire \M_target_pcb[10]~q ;
wire \A_pipe_flush_waddr_nxt~8_combout ;
wire \A_pipe_flush_waddr[8]~q ;
wire \D_pc_plus_one[8]~q ;
wire \E_extra_pc[8]~q ;
wire \M_pipe_flush_waddr[8]~q ;
wire \F_ic_tag_rd_addr_nxt[5]~15_combout ;
wire \F_pc[8]~q ;
wire \Add3~34 ;
wire \Add3~41_sumout ;
wire \Add0~30 ;
wire \Add0~25_sumout ;
wire \D_br_taken_waddr_partial[9]~q ;
wire \F_pc_nxt[9]~2_combout ;
wire \M_target_pcb[11]~q ;
wire \A_pipe_flush_waddr_nxt~10_combout ;
wire \A_pipe_flush_waddr[9]~q ;
wire \M_pipe_flush_waddr[9]~q ;
wire \F_pc_nxt[9]~3_combout ;
wire \F_pc[9]~q ;
wire \Add3~42 ;
wire \Add3~45_sumout ;
wire \D_pc_plus_one[10]~q ;
wire \Add0~26 ;
wire \Add0~41_sumout ;
wire \D_br_taken_waddr_partial[10]~q ;
wire \Add1~22_cout ;
wire \Add1~9_sumout ;
wire \F_pc_nxt[10]~4_combout ;
wire \M_target_pcb[12]~q ;
wire \A_pipe_flush_waddr_nxt~11_combout ;
wire \A_pipe_flush_waddr[10]~q ;
wire \M_pipe_flush_waddr[10]~q ;
wire \F_pc_nxt[10]~5_combout ;
wire \F_pc[10]~q ;
wire \Add3~46 ;
wire \Add3~49_sumout ;
wire \D_pc_plus_one[11]~q ;
wire \Add1~10 ;
wire \Add1~13_sumout ;
wire \F_pc_nxt[11]~6_combout ;
wire \M_target_pcb[13]~q ;
wire \A_pipe_flush_waddr_nxt~12_combout ;
wire \A_pipe_flush_waddr[11]~q ;
wire \M_pipe_flush_waddr[11]~q ;
wire \F_pc_nxt[11]~7_combout ;
wire \F_pc[11]~q ;
wire \Add3~50 ;
wire \Add3~53_sumout ;
wire \D_pc_plus_one[12]~q ;
wire \Add1~14 ;
wire \Add1~17_sumout ;
wire \F_pc_nxt[12]~8_combout ;
wire \Add7~53_sumout ;
wire \M_pc_plus_one[12]~q ;
wire \M_target_pcb[14]~q ;
wire \A_pipe_flush_waddr_nxt~13_combout ;
wire \A_pipe_flush_waddr[12]~q ;
wire \E_extra_pc[12]~q ;
wire \M_pipe_flush_waddr[12]~q ;
wire \F_pc_nxt[12]~9_combout ;
wire \F_pc[12]~q ;
wire \Add3~54 ;
wire \Add3~57_sumout ;
wire \D_pc_plus_one[13]~q ;
wire \Add1~18 ;
wire \Add1~5_sumout ;
wire \F_pc_nxt[13]~10_combout ;
wire \M_target_pcb[15]~q ;
wire \A_pipe_flush_waddr_nxt~14_combout ;
wire \A_pipe_flush_waddr[13]~q ;
wire \M_pipe_flush_waddr[13]~0_combout ;
wire \M_pipe_flush_waddr[13]~q ;
wire \F_pc_nxt[13]~11_combout ;
wire \F_pc[13]~q ;
wire \Add3~58 ;
wire \Add3~37_sumout ;
wire \D_pc_plus_one[14]~q ;
wire \Add1~6 ;
wire \Add1~1_sumout ;
wire \F_pc_nxt[14]~0_combout ;
wire \M_target_pcb[16]~q ;
wire \A_pipe_flush_waddr_nxt~9_combout ;
wire \A_pipe_flush_waddr[14]~q ;
wire \M_pipe_flush_waddr[14]~q ;
wire \F_pc_nxt[14]~1_combout ;
wire \F_pc[14]~q ;
wire \F_ic_hit~0_combout ;
wire \F_ic_hit~1_combout ;
wire \F_ic_hit~combout ;
wire \D_iw_valid~q ;
wire \F_kill~0_combout ;
wire \F_kill~combout ;
wire \F_issue~combout ;
wire \D_issue~q ;
wire \F_ic_tag_rd_addr_nxt[3]~0_combout ;
wire \F_ic_tag_rd_addr_nxt[0]~4_combout ;
wire \Add7~9_sumout ;
wire \M_pc_plus_one[3]~q ;
wire \M_target_pcb[5]~q ;
wire \A_pipe_flush_waddr_nxt~3_combout ;
wire \A_pipe_flush_waddr[3]~q ;
wire \M_pipe_flush_waddr[3]~q ;
wire \F_ic_tag_rd_addr_nxt[0]~5_combout ;
wire \F_pc[3]~q ;
wire \Add3~13_sumout ;
wire \Add0~13_sumout ;
wire \D_br_taken_waddr_partial[3]~q ;
wire \D_pc_plus_one[3]~q ;
wire \E_extra_pc[3]~q ;
wire \E_alu_result[5]~combout ;
wire \M_alu_result[5]~q ;
wire \D_src1_reg[5]~17_combout ;
wire \E_src1[5]~q ;
wire \E_rot_step1[5]~14_combout ;
wire \M_rot_prestep2[5]~q ;
wire \M_rot[5]~5_combout ;
wire \A_shift_rot_result~5_combout ;
wire \A_shift_rot_result[5]~q ;
wire \A_inst_result[5]~q ;
wire \A_mul_cell_p1[5]~q ;
wire \A_wr_data_unfiltered[5]~7_combout ;
wire \W_wr_data[5]~q ;
wire \D_src2_reg[5]~20_combout ;
wire \D_src2_reg[5]~21_combout ;
wire \E_src2[5]~q ;
wire \Add9~6 ;
wire \Add9~50 ;
wire \Add9~45_sumout ;
wire \E_alu_result~6_combout ;
wire \E_alu_result[7]~combout ;
wire \M_alu_result[7]~q ;
wire \D_src1_reg[7]~8_combout ;
wire \E_src1[7]~q ;
wire \E_rot_step1[7]~30_combout ;
wire \M_rot_prestep2[7]~q ;
wire \M_rot[7]~7_combout ;
wire \A_shift_rot_result~7_combout ;
wire \A_shift_rot_result[7]~q ;
wire \A_inst_result[7]~q ;
wire \A_mul_cell_p1[7]~q ;
wire \A_wr_data_unfiltered[7]~9_combout ;
wire \W_wr_data[7]~q ;
wire \D_src2_reg[7]~24_combout ;
wire \D_src2_reg[7]~25_combout ;
wire \E_src2[7]~q ;
wire \Equal316~3_combout ;
wire \Equal316~4_combout ;
wire \Equal316~5_combout ;
wire \Equal316~6_combout ;
wire \Equal316~7_combout ;
wire \Equal316~8_combout ;
wire \Equal316~9_combout ;
wire \Equal316~10_combout ;
wire \Equal316~11_combout ;
wire \Equal316~12_combout ;
wire \Equal316~13_combout ;
wire \Equal316~14_combout ;
wire \Equal316~15_combout ;
wire \E_compare_op[1]~q ;
wire \E_br_result~0_combout ;
wire \E_br_result~1_combout ;
wire \E_logic_result[0]~6_combout ;
wire \E_alu_result[0]~1_combout ;
wire \E_alu_result[0]~combout ;
wire \M_alu_result[0]~q ;
wire \D_src1_reg[0]~4_combout ;
wire \E_src1[0]~q ;
wire \E_rot_step1[2]~17_combout ;
wire \M_rot_prestep2[6]~q ;
wire \E_rot_step1[26]~19_combout ;
wire \M_rot_prestep2[30]~q ;
wire \M_rot[6]~6_combout ;
wire \A_shift_rot_result~6_combout ;
wire \A_shift_rot_result[6]~q ;
wire \A_inst_result[6]~q ;
wire \A_mul_cell_p1[6]~q ;
wire \A_wr_data_unfiltered[6]~8_combout ;
wire \W_wr_data[6]~q ;
wire \D_src2_reg[6]~22_combout ;
wire \D_src2_reg[6]~23_combout ;
wire \E_src2[6]~q ;
wire \Add9~49_sumout ;
wire \E_alu_result~5_combout ;
wire \E_alu_result[6]~combout ;
wire \M_alu_result[6]~q ;
wire \D_src1_reg[6]~18_combout ;
wire \E_src1[6]~q ;
wire \E_rot_step1[6]~22_combout ;
wire \M_rot_prestep2[10]~q ;
wire \E_rot_step1[22]~18_combout ;
wire \M_rot_prestep2[26]~q ;
wire \M_rot[2]~16_combout ;
wire \A_shift_rot_result~16_combout ;
wire \A_shift_rot_result[10]~q ;
wire \A_inst_result[10]~q ;
wire \A_mul_cell_p1[10]~q ;
wire \A_wr_data_unfiltered[10]~18_combout ;
wire \W_wr_data[10]~q ;
wire \D_src2_reg[10]~43_combout ;
wire \D_src2_reg[10]~44_combout ;
wire \E_src2[10]~q ;
wire \Add9~37_sumout ;
wire \E_alu_result~13_combout ;
wire \E_alu_result[10]~combout ;
wire \M_alu_result[10]~q ;
wire \D_src1_reg[10]~12_combout ;
wire \E_src1[10]~q ;
wire \E_rot_step1[10]~23_combout ;
wire \M_rot_prestep2[14]~q ;
wire \M_rot[6]~30_combout ;
wire \A_shift_rot_result~30_combout ;
wire \A_shift_rot_result[14]~q ;
wire \A_inst_result[14]~q ;
wire \A_mul_cell_p1[14]~q ;
wire \A_wr_data_unfiltered[14]~32_combout ;
wire \W_wr_data[14]~q ;
wire \D_src2_reg[14]~68_combout ;
wire \D_src2_reg[14]~69_combout ;
wire \E_src2[14]~q ;
wire \Add9~21_sumout ;
wire \E_alu_result~23_combout ;
wire \E_alu_result[14]~combout ;
wire \M_alu_result[14]~q ;
wire \D_src1_reg[14]~30_combout ;
wire \E_src1[14]~q ;
wire \E_rot_step1[14]~20_combout ;
wire \M_rot_prestep2[18]~q ;
wire \M_rot[2]~25_combout ;
wire \A_shift_rot_result~25_combout ;
wire \A_shift_rot_result[18]~q ;
wire \A_inst_result[18]~q ;
wire \Add12~53_sumout ;
wire \A_wr_data_unfiltered[18]~27_combout ;
wire \W_wr_data[18]~q ;
wire \D_src2_reg[18]~60_combout ;
wire \Add9~125_sumout ;
wire \D_src2[18]~35_combout ;
wire \D_src2[18]~36_combout ;
wire \D_src2[18]~25_combout ;
wire \E_src2[18]~q ;
wire \E_logic_result[18]~11_combout ;
wire \E_alu_result[18]~combout ;
wire \M_alu_result[18]~q ;
wire \D_src1_reg[18]~25_combout ;
wire \E_src1[18]~q ;
wire \E_rot_step1[18]~21_combout ;
wire \M_rot_prestep2[22]~q ;
wire \M_rot[6]~8_combout ;
wire \A_shift_rot_result~8_combout ;
wire \A_shift_rot_result[22]~q ;
wire \A_inst_result[22]~q ;
wire \Add11~22 ;
wire \Add11~1_sumout ;
wire \A_mul_s1[6]~q ;
wire \A_mul_cell_p3[6]~q ;
wire \Add12~22 ;
wire \Add12~1_sumout ;
wire \A_wr_data_unfiltered[22]~10_combout ;
wire \W_wr_data[22]~q ;
wire \D_src1_reg[22]~1_combout ;
wire \E_src1[22]~q ;
wire \E_logic_result[22]~1_combout ;
wire \Add9~94 ;
wire \Add9~77_sumout ;
wire \E_alu_result[22]~combout ;
wire \M_alu_result[22]~q ;
wire \D_src2_reg[22]~26_combout ;
wire \D_src2[22]~41_combout ;
wire \D_src2[22]~42_combout ;
wire \D_src2[22]~1_combout ;
wire \E_src2[22]~q ;
wire \Add9~78 ;
wire \Add9~81_sumout ;
wire \E_alu_result[23]~combout ;
wire \M_alu_result[23]~q ;
wire \A_slow_inst_result_nxt[23]~36_combout ;
wire \A_slow_inst_result_nxt[23]~9_combout ;
wire \A_slow_inst_result[23]~q ;
wire \M_rot[7]~9_combout ;
wire \A_shift_rot_result~9_combout ;
wire \A_shift_rot_result[23]~q ;
wire \A_inst_result[23]~q ;
wire \Add11~2 ;
wire \Add11~5_sumout ;
wire \A_mul_s1[7]~q ;
wire \A_mul_cell_p3[7]~q ;
wire \Add12~2 ;
wire \Add12~5_sumout ;
wire \A_wr_data_unfiltered[23]~11_combout ;
wire \W_wr_data[23]~q ;
wire \D_src1_reg[23]~2_combout ;
wire \E_src1[23]~q ;
wire \E_logic_result[23]~2_combout ;
wire \E_alu_result~7_combout ;
wire \D_src2_reg[23]~27_combout ;
wire \D_src2_reg[0]~9_combout ;
wire \D_src2_reg[23]~28_combout ;
wire \D_src2[23]~2_combout ;
wire \D_src2[23]~3_combout ;
wire \E_src2[23]~q ;
wire \Add9~82 ;
wire \Add9~85_sumout ;
wire \E_alu_result[24]~combout ;
wire \M_alu_result[24]~q ;
wire \A_slow_inst_result_nxt[24]~37_combout ;
wire \A_slow_inst_result_nxt[24]~10_combout ;
wire \A_slow_inst_result[24]~q ;
wire \E_rot_pass3~0_combout ;
wire \M_rot_pass3~q ;
wire \E_rot_sel_fill3~0_combout ;
wire \M_rot_sel_fill3~q ;
wire \M_rot[0]~10_combout ;
wire \A_shift_rot_result~10_combout ;
wire \A_shift_rot_result[24]~q ;
wire \A_inst_result[24]~q ;
wire \Add11~6 ;
wire \Add11~9_sumout ;
wire \A_mul_s1[8]~q ;
wire \A_mul_cell_p3[8]~q ;
wire \Add12~6 ;
wire \Add12~9_sumout ;
wire \A_wr_data_unfiltered[24]~12_combout ;
wire \W_wr_data[24]~q ;
wire \D_src1_reg[24]~3_combout ;
wire \E_src1[24]~q ;
wire \E_logic_result[24]~3_combout ;
wire \E_alu_result~8_combout ;
wire \D_src2_reg[24]~29_combout ;
wire \D_src2_reg[24]~30_combout ;
wire \D_src2[24]~4_combout ;
wire \D_src2[24]~5_combout ;
wire \E_src2[24]~q ;
wire \Add9~86 ;
wire \Add9~89_sumout ;
wire \E_alu_result[25]~combout ;
wire \M_alu_result[25]~q ;
wire \A_slow_inst_result_nxt[25]~39_combout ;
wire \A_slow_inst_result_nxt[25]~11_combout ;
wire \A_slow_inst_result[25]~q ;
wire \M_rot[1]~11_combout ;
wire \A_shift_rot_result~11_combout ;
wire \A_shift_rot_result[25]~q ;
wire \A_inst_result[25]~q ;
wire \Add11~10 ;
wire \Add11~13_sumout ;
wire \A_mul_s1[9]~q ;
wire \A_mul_cell_p3[9]~q ;
wire \Add12~10 ;
wire \Add12~13_sumout ;
wire \A_wr_data_unfiltered[25]~13_combout ;
wire \W_wr_data[25]~q ;
wire \D_src1_reg[25]~5_combout ;
wire \E_src1[25]~q ;
wire \E_alu_result~9_combout ;
wire \D_src2_reg[25]~31_combout ;
wire \D_src2_reg[25]~32_combout ;
wire \D_src2[25]~6_combout ;
wire \D_src2[25]~7_combout ;
wire \E_src2[25]~q ;
wire \Add9~90 ;
wire \Add9~105_sumout ;
wire \E_alu_result[26]~combout ;
wire \M_alu_result[26]~q ;
wire \A_slow_inst_result_nxt[26]~24_combout ;
wire \A_slow_inst_result_nxt[26]~16_combout ;
wire \A_slow_inst_result[26]~q ;
wire \M_rot[2]~20_combout ;
wire \A_shift_rot_result~20_combout ;
wire \A_shift_rot_result[26]~q ;
wire \A_inst_result[26]~q ;
wire \Add11~14 ;
wire \Add11~33_sumout ;
wire \A_mul_s1[10]~q ;
wire \A_mul_cell_p3[10]~q ;
wire \Add12~14 ;
wire \Add12~33_sumout ;
wire \A_wr_data_unfiltered[26]~22_combout ;
wire \W_wr_data[26]~q ;
wire \D_src1_reg[26]~19_combout ;
wire \E_src1[26]~q ;
wire \E_alu_result~17_combout ;
wire \D_src2_reg[26]~52_combout ;
wire \D_src2_reg[26]~53_combout ;
wire \D_src2[26]~17_combout ;
wire \D_src2[26]~18_combout ;
wire \E_src2[26]~q ;
wire \Add9~106 ;
wire \Add9~101_sumout ;
wire \E_alu_result[27]~combout ;
wire \M_alu_result[27]~q ;
wire \A_slow_inst_result_nxt[27]~25_combout ;
wire \A_slow_inst_result_nxt[27]~15_combout ;
wire \A_slow_inst_result[27]~q ;
wire \M_rot[3]~17_combout ;
wire \A_shift_rot_result~17_combout ;
wire \A_shift_rot_result[27]~q ;
wire \A_inst_result[27]~q ;
wire \Add11~34 ;
wire \Add11~29_sumout ;
wire \A_mul_s1[11]~q ;
wire \A_mul_cell_p3[11]~q ;
wire \Add12~34 ;
wire \Add12~29_sumout ;
wire \A_wr_data_unfiltered[27]~19_combout ;
wire \W_wr_data[27]~q ;
wire \D_src1_reg[27]~13_combout ;
wire \E_src1[27]~q ;
wire \E_alu_result~14_combout ;
wire \D_src2_reg[27]~45_combout ;
wire \D_src2_reg[27]~34_combout ;
wire \D_src2_reg[27]~46_combout ;
wire \D_src2_reg[27]~47_combout ;
wire \D_src2[27]~14_combout ;
wire \D_src2[27]~15_combout ;
wire \E_src2[27]~q ;
wire \Add9~102 ;
wire \Add9~97_sumout ;
wire \E_alu_result[28]~combout ;
wire \M_alu_result[28]~q ;
wire \A_slow_inst_result_nxt[28]~26_combout ;
wire \A_slow_inst_result_nxt[28]~14_combout ;
wire \A_slow_inst_result[28]~q ;
wire \M_rot[4]~15_combout ;
wire \A_shift_rot_result~15_combout ;
wire \A_shift_rot_result[28]~q ;
wire \A_inst_result[28]~q ;
wire \Add11~30 ;
wire \Add11~25_sumout ;
wire \A_mul_s1[12]~q ;
wire \A_mul_cell_p3[12]~q ;
wire \Add12~30 ;
wire \Add12~25_sumout ;
wire \A_wr_data_unfiltered[28]~17_combout ;
wire \W_wr_data[28]~q ;
wire \D_src1_reg[28]~11_combout ;
wire \E_src1[28]~q ;
wire \E_alu_result~12_combout ;
wire \D_src2_reg[28]~40_combout ;
wire \D_src2_reg[28]~41_combout ;
wire \D_src2_reg[28]~42_combout ;
wire \D_src2[28]~12_combout ;
wire \D_src2[28]~13_combout ;
wire \E_src2[28]~q ;
wire \Add9~98 ;
wire \Add9~129_sumout ;
wire \E_alu_result[29]~combout ;
wire \M_alu_result[29]~q ;
wire \A_slow_inst_result_nxt[29]~28_combout ;
wire \A_slow_inst_result_nxt[29]~23_combout ;
wire \A_slow_inst_result[29]~q ;
wire \M_rot[5]~31_combout ;
wire \A_shift_rot_result~31_combout ;
wire \A_shift_rot_result[29]~q ;
wire \A_inst_result[29]~q ;
wire \Add11~26 ;
wire \Add11~61_sumout ;
wire \A_mul_s1[13]~q ;
wire \A_mul_cell_p3[13]~q ;
wire \Add12~26 ;
wire \Add12~61_sumout ;
wire \A_wr_data_unfiltered[29]~33_combout ;
wire \W_wr_data[29]~q ;
wire \D_src1_reg[29]~31_combout ;
wire \E_src1[29]~q ;
wire \E_alu_result~24_combout ;
wire \D_src2_reg[29]~70_combout ;
wire \D_src2_reg[29]~71_combout ;
wire \D_src2_reg[29]~72_combout ;
wire \D_src2[29]~27_combout ;
wire \D_src2[29]~28_combout ;
wire \E_src2[29]~q ;
wire \Add9~130 ;
wire \Add9~121_sumout ;
wire \D_src2_reg[30]~57_combout ;
wire \A_slow_inst_result_nxt[30]~31_combout ;
wire \A_slow_inst_result_nxt[30]~20_combout ;
wire \A_slow_inst_result[30]~q ;
wire \M_rot[6]~24_combout ;
wire \A_shift_rot_result~24_combout ;
wire \A_shift_rot_result[30]~q ;
wire \A_inst_result[30]~q ;
wire \Add11~62 ;
wire \Add11~49_sumout ;
wire \A_mul_s1[14]~q ;
wire \A_mul_cell_p3[14]~q ;
wire \Add12~62 ;
wire \Add12~49_sumout ;
wire \A_wr_data_unfiltered[30]~26_combout ;
wire \W_wr_data[30]~q ;
wire \D_src2_reg[30]~58_combout ;
wire \D_src2_reg[30]~59_combout ;
wire \D_src2[30]~22_combout ;
wire \D_src2[30]~23_combout ;
wire \E_src2[30]~q ;
wire \E_logic_result[30]~5_combout ;
wire \E_alu_result~18_combout ;
wire \E_alu_result[30]~combout ;
wire \M_alu_result[30]~q ;
wire \D_src1_reg[30]~23_combout ;
wire \E_src1[30]~q ;
wire \E_rot_step1[30]~16_combout ;
wire \M_rot_prestep2[2]~q ;
wire \M_rot[2]~2_combout ;
wire \A_shift_rot_result~2_combout ;
wire \A_shift_rot_result[2]~q ;
wire \Equal327~0_combout ;
wire \latched_oci_tb_hbreak_req_next~0_combout ;
wire \latched_oci_tb_hbreak_req~q ;
wire \A_exc_norm_intr_pri5_nxt~0_combout ;
wire \A_exc_norm_intr_pri5~q ;
wire \A_exc_trap_inst_pri15_nxt~0_combout ;
wire \A_exc_trap_inst_pri15~q ;
wire \A_exc_illegal_inst_pri15_nxt~0_combout ;
wire \A_exc_illegal_inst_pri15~q ;
wire \A_exc_highest_pri_cause_code[0]~0_combout ;
wire \A_exc_active_no_break~combout ;
wire \W_exception_reg_cause[0]~q ;
wire \E_control_reg_rddata_muxed[2]~2_combout ;
wire \M_control_reg_rddata[2]~q ;
wire \M_inst_result[2]~2_combout ;
wire \A_inst_result[2]~q ;
wire \A_mul_cell_p1[2]~q ;
wire \A_wr_data_unfiltered[2]~4_combout ;
wire \W_wr_data[2]~q ;
wire \D_src1_reg[2]~6_combout ;
wire \E_src1[2]~q ;
wire \Add9~57_sumout ;
wire \E_alu_result~2_combout ;
wire \E_alu_result[2]~combout ;
wire \D_src2_reg[2]~14_combout ;
wire \D_src2[2]~46_combout ;
wire \D_src2[2]~8_combout ;
wire \E_src2[2]~q ;
wire \E_rot_mask[4]~4_combout ;
wire \M_rot_mask[4]~q ;
wire \M_rot[4]~4_combout ;
wire \A_shift_rot_result~4_combout ;
wire \A_shift_rot_result[4]~q ;
wire \A_exc_highest_pri_cause_code[1]~1_combout ;
wire \W_exception_reg_cause[2]~0_combout ;
wire \W_exception_reg_cause[2]~q ;
wire \E_control_reg_rddata_muxed[4]~4_combout ;
wire \M_control_reg_rddata[4]~q ;
wire \M_inst_result[4]~4_combout ;
wire \A_inst_result[4]~q ;
wire \A_mul_cell_p1[4]~q ;
wire \A_wr_data_unfiltered[4]~6_combout ;
wire \W_wr_data[4]~q ;
wire \D_src1_reg[4]~16_combout ;
wire \E_src1[4]~q ;
wire \Add9~1_sumout ;
wire \E_alu_result~3_combout ;
wire \E_alu_result[4]~combout ;
wire \D_src2_reg[4]~18_combout ;
wire \D_src2[4]~43_combout ;
wire \D_src2[4]~16_combout ;
wire \E_src2[4]~q ;
wire \E_rot_sel_fill0~0_combout ;
wire \M_rot_sel_fill0~q ;
wire \M_rot[3]~3_combout ;
wire \A_shift_rot_result~3_combout ;
wire \A_shift_rot_result[3]~q ;
wire \W_exception_reg_cause[1]~q ;
wire \E_control_reg_rddata_muxed[3]~3_combout ;
wire \M_control_reg_rddata[3]~q ;
wire \M_inst_result[3]~3_combout ;
wire \A_inst_result[3]~q ;
wire \A_mul_cell_p1[3]~q ;
wire \A_wr_data_unfiltered[3]~5_combout ;
wire \W_wr_data[3]~q ;
wire \D_src1_reg[3]~0_combout ;
wire \E_src1[3]~q ;
wire \Add9~53_sumout ;
wire \E_alu_result[3]~combout ;
wire \D_src2_reg[3]~16_combout ;
wire \D_src2[3]~45_combout ;
wire \D_src2[3]~0_combout ;
wire \E_src2[3]~q ;
wire \E_rot_pass0~0_combout ;
wire \M_rot_pass0~q ;
wire \M_rot[0]~0_combout ;
wire \A_shift_rot_result~0_combout ;
wire \A_shift_rot_result[0]~q ;
wire \W_estatus_reg_pie_nxt~0_combout ;
wire \W_estatus_reg_pie_nxt~1_combout ;
wire \W_estatus_reg_pie~q ;
wire \W_bstatus_reg_pie_nxt~0_combout ;
wire \W_bstatus_reg_pie_nxt~1_combout ;
wire \W_bstatus_reg_pie~q ;
wire \D_control_reg_rddata_muxed[0]~0_combout ;
wire \D_control_reg_rddata_muxed[0]~1_combout ;
wire \E_control_reg_rddata[0]~q ;
wire \E_control_reg_rddata_muxed[0]~0_combout ;
wire \M_control_reg_rddata[0]~q ;
wire \M_inst_result[0]~0_combout ;
wire \A_inst_result[0]~q ;
wire \A_mul_cell_p1[0]~q ;
wire \A_wr_data_unfiltered[0]~2_combout ;
wire \W_wr_data[0]~q ;
wire \D_src2_reg[0]~10_combout ;
wire \D_src2[0]~47_combout ;
wire \E_src2[0]~q ;
wire \Add9~65_sumout ;
wire \M_mem_baddr[0]~q ;
wire \M_ld_align_sh8~combout ;
wire \A_ld_align_sh8~q ;
wire \A_slow_inst_result_nxt[1]~1_combout ;
wire \A_slow_inst_result[1]~q ;
wire \M_rot[1]~1_combout ;
wire \A_shift_rot_result~1_combout ;
wire \A_shift_rot_result[1]~q ;
wire \W_ienable_reg_irq1~q ;
wire \W_ipending_reg_irq1_nxt~combout ;
wire \W_ipending_reg_irq1~q ;
wire \D_control_reg_rddata_muxed[1]~2_combout ;
wire \E_control_reg_rddata[1]~q ;
wire \E_control_reg_rddata_muxed[1]~1_combout ;
wire \M_control_reg_rddata[1]~q ;
wire \M_inst_result[1]~1_combout ;
wire \A_inst_result[1]~q ;
wire \A_mul_cell_p1[1]~q ;
wire \A_wr_data_unfiltered[1]~3_combout ;
wire \W_wr_data[1]~q ;
wire \D_src1_reg[1]~24_combout ;
wire \E_src1[1]~q ;
wire \E_logic_result[1]~7_combout ;
wire \E_alu_result[1]~combout ;
wire \D_src2_reg[1]~12_combout ;
wire \D_src2[1]~44_combout ;
wire \D_src2[1]~24_combout ;
wire \E_src2[1]~q ;
wire \Add9~69_sumout ;
wire \M_mem_baddr[1]~q ;
wire \A_mem_baddr[1]~q ;
wire \A_mem_baddr[0]~q ;
wire \A_ctrl_ld16~q ;
wire \A_slow_ld_data_sign_bit~0_combout ;
wire \M_ctrl_ld_signed~q ;
wire \A_ctrl_ld_signed~q ;
wire \A_slow_ld_data_fill_bit~0_combout ;
wire \A_slow_inst_result_nxt[31]~38_combout ;
wire \A_slow_inst_result_nxt[31]~12_combout ;
wire \A_slow_inst_result[31]~q ;
wire \M_rot[7]~12_combout ;
wire \A_shift_rot_result~12_combout ;
wire \A_shift_rot_result[31]~q ;
wire \A_inst_result[31]~q ;
wire \Add11~50 ;
wire \Add11~17_sumout ;
wire \A_mul_s1[15]~q ;
wire \A_mul_cell_p3[15]~q ;
wire \Add12~50 ;
wire \Add12~17_sumout ;
wire \A_wr_data_unfiltered[31]~14_combout ;
wire \W_wr_data[31]~q ;
wire \D_src1_reg[31]~7_combout ;
wire \E_src1[31]~q ;
wire \Add9~122 ;
wire \Add9~73_sumout ;
wire \D_src2_reg[31]~33_combout ;
wire \D_src2_reg[31]~35_combout ;
wire \D_src2_reg[31]~36_combout ;
wire \D_src2[31]~9_combout ;
wire \D_src2[31]~10_combout ;
wire \E_src2[31]~q ;
wire \Add9~74 ;
wire \Add9~61_sumout ;
wire \E_bht_data[1]~q ;
wire \E_ctrl_br_cond~q ;
wire \E_br_mispredict~0_combout ;
wire \M_pipe_flush_nxt~combout ;
wire \M_pipe_flush~q ;
wire \D_ctrl_shift_rot~1_combout ;
wire \D_ctrl_late_result~1_combout ;
wire \D_ctrl_late_result~0_combout ;
wire \E_ctrl_late_result~q ;
wire \D_data_depend~0_combout ;
wire \M_ctrl_late_result~q ;
wire \D_data_depend~1_combout ;
wire \D_valid~combout ;
wire \E_valid_from_D~q ;
wire \E_valid~combout ;
wire \M_valid_from_E~q ;
wire \M_exc_allowed~0_combout ;
wire \A_exc_allowed~q ;
wire \wait_for_one_post_bret_inst~1_combout ;
wire \wait_for_one_post_bret_inst~q ;
wire \wait_for_one_post_bret_inst~0_combout ;
wire \hbreak_req~0_combout ;
wire \M_exc_any~combout ;
wire \A_exc_any~q ;
wire \M_iw[11]~q ;
wire \A_iw[11]~q ;
wire \M_iw[5]~q ;
wire \A_iw[5]~q ;
wire \M_iw[0]~q ;
wire \A_iw[0]~q ;
wire \M_iw[16]~q ;
wire \A_iw[16]~q ;
wire \M_iw[15]~q ;
wire \A_iw[15]~q ;
wire \M_iw[13]~q ;
wire \A_iw[13]~q ;
wire \M_iw[12]~q ;
wire \A_iw[12]~q ;
wire \A_op_eret~0_combout ;
wire \M_iw[4]~q ;
wire \A_iw[4]~q ;
wire \M_iw[3]~q ;
wire \A_iw[3]~q ;
wire \M_iw[2]~q ;
wire \A_iw[2]~q ;
wire \M_iw[1]~q ;
wire \A_iw[1]~q ;
wire \A_op_eret~1_combout ;
wire \A_op_eret~2_combout ;
wire \W_status_reg_pie_nxt~0_combout ;
wire \M_iw[14]~q ;
wire \A_iw[14]~q ;
wire \W_status_reg_pie_nxt~1_combout ;
wire \W_status_reg_pie_nxt~2_combout ;
wire \W_status_reg_pie_nxt~3_combout ;
wire \W_status_reg_pie~q ;
wire \norm_intr_req~0_combout ;
wire \M_norm_intr_req~q ;
wire \M_valid~0_combout ;
wire \M_data_master_start_stall~0_combout ;
wire \E_ctrl_ld_st~0_combout ;
wire \M_ctrl_ld_st~q ;
wire \E_ctrl_st~0_combout ;
wire \M_ctrl_st~q ;
wire \A_ctrl_st~q ;
wire \M_data_master_start_stall~combout ;
wire \A_data_master_started_stall~q ;
wire \av_ld_data_transfer~0_combout ;
wire \av_ld_aligning_data~q ;
wire \A_mem_stall_nxt~0_combout ;
wire \A_mem_stall_nxt~1_combout ;
wire \A_mem_stall~q ;
wire \F_stall~0_combout ;
wire \D_iw[5]~q ;
wire \D_ctrl_cmp~0_combout ;
wire \D_ctrl_cmp~1_combout ;
wire \D_ctrl_cmp~3_combout ;
wire \D_ctrl_cmp~2_combout ;
wire \E_ctrl_cmp~q ;
wire \D_src2_reg[0]~3_combout ;
wire \D_src2_reg[0]~11_combout ;
wire \E_src2_reg[0]~q ;
wire \M_st_data[0]~q ;
wire \M_mem_baddr[4]~q ;
wire \M_mem_baddr[5]~q ;
wire \M_mem_baddr[8]~q ;
wire \M_mem_baddr[16]~q ;
wire \M_mem_baddr[15]~q ;
wire \M_mem_baddr[14]~q ;
wire \M_mem_baddr[13]~q ;
wire \M_mem_baddr[12]~q ;
wire \M_mem_baddr[11]~q ;
wire \M_mem_baddr[10]~q ;
wire \M_mem_baddr[9]~q ;
wire \M_mem_baddr[7]~q ;
wire \M_mem_baddr[6]~q ;
wire \d_write_nxt~combout ;
wire \M_mem_baddr[3]~q ;
wire \M_mem_baddr[2]~q ;
wire \D_src2_reg[1]~13_combout ;
wire \E_src2_reg[1]~q ;
wire \M_st_data[1]~q ;
wire \D_src2_reg[2]~15_combout ;
wire \E_src2_reg[2]~q ;
wire \M_st_data[2]~q ;
wire \D_src2_reg[3]~17_combout ;
wire \E_src2_reg[3]~q ;
wire \M_st_data[3]~q ;
wire \D_src2_reg[4]~19_combout ;
wire \E_src2_reg[4]~q ;
wire \M_st_data[4]~q ;
wire \E_src2_reg[5]~q ;
wire \M_st_data[5]~q ;
wire \E_src2_reg[6]~q ;
wire \M_st_data[6]~q ;
wire \E_src2_reg[7]~q ;
wire \M_st_data[7]~q ;
wire \d_read_nxt~combout ;
wire \W_debug_mode_nxt~0_combout ;
wire \F_ic_fill_same_tag_line~0_combout ;
wire \F_ic_fill_same_tag_line~1_combout ;
wire \F_ic_fill_same_tag_line~2_combout ;
wire \F_ic_fill_same_tag_line~3_combout ;
wire \F_ic_fill_same_tag_line~4_combout ;
wire \F_ic_fill_same_tag_line~5_combout ;
wire \F_ic_fill_same_tag_line~combout ;
wire \D_ic_fill_same_tag_line~q ;
wire \E_ctrl_invalidate_i~0_combout ;
wire \E_ctrl_invalidate_i~1_combout ;
wire \M_ctrl_invalidate_i~q ;
wire \A_ctrl_invalidate_i~q ;
wire \ic_fill_prevent_refill_nxt~combout ;
wire \ic_fill_prevent_refill~q ;
wire \D_ic_fill_starting~0_combout ;
wire \D_ic_fill_starting~combout ;
wire \ic_fill_initial_offset[2]~q ;
wire \D_ic_fill_starting_d1~q ;
wire \ic_fill_initial_offset[0]~q ;
wire \ic_fill_dp_offset_nxt[0]~1_combout ;
wire \i_readdatavalid_d1~q ;
wire \ic_fill_dp_offset_en~0_combout ;
wire \ic_fill_dp_offset[0]~q ;
wire \ic_fill_initial_offset[1]~q ;
wire \ic_fill_dp_offset_nxt[1]~2_combout ;
wire \ic_fill_dp_offset[1]~q ;
wire \ic_fill_dp_offset[2]~q ;
wire \ic_fill_dp_offset_nxt[2]~0_combout ;
wire \ic_fill_active_nxt~0_combout ;
wire \ic_fill_active_nxt~1_combout ;
wire \ic_fill_active~q ;
wire \ic_fill_ap_cnt_nxt[0]~3_combout ;
wire \ic_fill_ap_offset[2]~0_combout ;
wire \ic_fill_ap_cnt[0]~q ;
wire \ic_fill_ap_cnt_nxt[1]~2_combout ;
wire \ic_fill_ap_cnt[1]~q ;
wire \ic_fill_ap_cnt_nxt[2]~1_combout ;
wire \ic_fill_ap_cnt[2]~q ;
wire \ic_fill_ap_cnt_nxt[3]~0_combout ;
wire \ic_fill_ap_cnt[3]~q ;
wire \i_read_nxt~0_combout ;
wire \i_read_nxt~1_combout ;
wire \ic_fill_ap_offset_nxt[0]~0_combout ;
wire \ic_tag_wraddress_nxt~0_combout ;
wire \ic_fill_ap_offset_nxt[2]~1_combout ;
wire \ic_fill_ap_offset_nxt[1]~2_combout ;
wire \ic_tag_wraddress_nxt~1_combout ;
wire \ic_tag_wraddress_nxt~2_combout ;
wire \ic_tag_wraddress_nxt~3_combout ;
wire \ic_tag_wraddress_nxt~4_combout ;
wire \ic_tag_wraddress_nxt~5_combout ;
wire \D_ctrl_mem16~0_combout ;
wire \E_ctrl_mem16~q ;
wire \D_ctrl_mem8~0_combout ;
wire \E_ctrl_mem8~q ;
wire \E_mem_byte_en~0_combout ;
wire \M_mem_byte_en[0]~q ;
wire \D_src2_reg[16]~73_combout ;
wire \E_src2_reg[16]~q ;
wire \E_st_data[23]~0_combout ;
wire \M_st_data[16]~q ;
wire \D_src2_reg[22]~74_combout ;
wire \E_src2_reg[22]~q ;
wire \M_st_data[22]~q ;
wire \E_mem_byte_en[2]~1_combout ;
wire \M_mem_byte_en[2]~q ;
wire \D_src2_reg[23]~75_combout ;
wire \E_src2_reg[23]~q ;
wire \M_st_data[23]~q ;
wire \E_src2_reg[8]~q ;
wire \D_src2_reg[24]~76_combout ;
wire \E_src2_reg[24]~q ;
wire \E_st_data[24]~1_combout ;
wire \M_st_data[24]~q ;
wire \E_mem_byte_en[3]~2_combout ;
wire \M_mem_byte_en[3]~q ;
wire \E_src2_reg[9]~q ;
wire \D_src2_reg[25]~77_combout ;
wire \E_src2_reg[25]~q ;
wire \E_st_data[25]~2_combout ;
wire \M_st_data[25]~q ;
wire \E_src2_reg[15]~q ;
wire \D_src2_reg[31]~89_combout ;
wire \D_src2_reg[31]~78_combout ;
wire \E_src2_reg[31]~q ;
wire \E_st_data[31]~3_combout ;
wire \M_st_data[31]~q ;
wire \D_src2_reg[21]~79_combout ;
wire \E_src2_reg[21]~q ;
wire \M_st_data[21]~q ;
wire \E_src2_reg[11]~q ;
wire \M_st_data[11]~q ;
wire \E_mem_byte_en[1]~3_combout ;
wire \M_mem_byte_en[1]~q ;
wire \E_src2_reg[12]~q ;
wire \D_src2_reg[28]~80_combout ;
wire \E_src2_reg[28]~q ;
wire \E_st_data[28]~4_combout ;
wire \M_st_data[28]~q ;
wire \E_src2_reg[10]~q ;
wire \M_st_data[10]~q ;
wire \D_src2_reg[27]~81_combout ;
wire \E_src2_reg[27]~q ;
wire \E_st_data[27]~5_combout ;
wire \M_st_data[27]~q ;
wire \M_st_data[8]~q ;
wire \M_st_data[9]~q ;
wire \D_src2_reg[26]~82_combout ;
wire \E_src2_reg[26]~q ;
wire \E_st_data[26]~6_combout ;
wire \M_st_data[26]~q ;
wire \D_src2_reg[20]~83_combout ;
wire \E_src2_reg[20]~q ;
wire \M_st_data[20]~q ;
wire \D_src2_reg[19]~84_combout ;
wire \E_src2_reg[19]~q ;
wire \M_st_data[19]~q ;
wire \D_src2_reg[17]~85_combout ;
wire \E_src2_reg[17]~q ;
wire \M_st_data[17]~q ;
wire \E_src2_reg[14]~q ;
wire \D_src2_reg[30]~86_combout ;
wire \E_src2_reg[30]~q ;
wire \E_st_data[30]~7_combout ;
wire \M_st_data[30]~q ;
wire \D_src2_reg[18]~87_combout ;
wire \E_src2_reg[18]~q ;
wire \M_st_data[18]~q ;
wire \M_st_data[15]~q ;
wire \M_st_data[12]~q ;
wire \E_src2_reg[13]~q ;
wire \M_st_data[13]~q ;
wire \M_st_data[14]~q ;
wire \D_src2_reg[29]~88_combout ;
wire \E_src2_reg[29]~q ;
wire \E_st_data[29]~8_combout ;
wire \M_st_data[29]~q ;


first_nios2_system_first_nios2_system_cpu_cpu_register_bank_a_module first_nios2_system_cpu_cpu_register_bank_a(
	.q_b_3(\first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[3] ),
	.q_b_22(\first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[22] ),
	.q_b_23(\first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[23] ),
	.q_b_24(\first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[24] ),
	.q_b_0(\first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[0] ),
	.q_b_25(\first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[25] ),
	.q_b_2(\first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[2] ),
	.q_b_31(\first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[31] ),
	.q_b_7(\first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[7] ),
	.q_b_21(\first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[21] ),
	.q_b_11(\first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[11] ),
	.q_b_28(\first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[28] ),
	.q_b_10(\first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[10] ),
	.q_b_27(\first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[27] ),
	.q_b_8(\first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[8] ),
	.q_b_9(\first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[9] ),
	.q_b_4(\first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[4] ),
	.q_b_5(\first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[5] ),
	.q_b_6(\first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[6] ),
	.q_b_26(\first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[26] ),
	.q_b_20(\first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[20] ),
	.q_b_19(\first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[19] ),
	.q_b_17(\first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[17] ),
	.q_b_30(\first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[30] ),
	.q_b_1(\first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[1] ),
	.q_b_18(\first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[18] ),
	.q_b_16(\first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[16] ),
	.q_b_15(\first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[15] ),
	.q_b_12(\first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[12] ),
	.q_b_13(\first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[13] ),
	.q_b_14(\first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[14] ),
	.q_b_29(\first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[29] ),
	.A_wr_data_unfiltered_0(\A_wr_data_unfiltered[0]~2_combout ),
	.A_wr_data_unfiltered_1(\A_wr_data_unfiltered[1]~3_combout ),
	.A_wr_data_unfiltered_2(\A_wr_data_unfiltered[2]~4_combout ),
	.A_wr_data_unfiltered_3(\A_wr_data_unfiltered[3]~5_combout ),
	.A_wr_data_unfiltered_4(\A_wr_data_unfiltered[4]~6_combout ),
	.A_wr_data_unfiltered_5(\A_wr_data_unfiltered[5]~7_combout ),
	.A_wr_data_unfiltered_6(\A_wr_data_unfiltered[6]~8_combout ),
	.A_wr_data_unfiltered_7(\A_wr_data_unfiltered[7]~9_combout ),
	.A_wr_data_unfiltered_22(\A_wr_data_unfiltered[22]~10_combout ),
	.A_wr_data_unfiltered_23(\A_wr_data_unfiltered[23]~11_combout ),
	.A_wr_data_unfiltered_24(\A_wr_data_unfiltered[24]~12_combout ),
	.A_wr_data_unfiltered_25(\A_wr_data_unfiltered[25]~13_combout ),
	.A_wr_data_unfiltered_31(\A_wr_data_unfiltered[31]~14_combout ),
	.A_wr_data_unfiltered_21(\A_wr_data_unfiltered[21]~15_combout ),
	.A_wr_data_unfiltered_11(\A_wr_data_unfiltered[11]~16_combout ),
	.A_wr_data_unfiltered_28(\A_wr_data_unfiltered[28]~17_combout ),
	.A_wr_data_unfiltered_10(\A_wr_data_unfiltered[10]~18_combout ),
	.A_wr_data_unfiltered_27(\A_wr_data_unfiltered[27]~19_combout ),
	.A_wr_data_unfiltered_8(\A_wr_data_unfiltered[8]~20_combout ),
	.A_wr_data_unfiltered_9(\A_wr_data_unfiltered[9]~21_combout ),
	.A_wr_data_unfiltered_26(\A_wr_data_unfiltered[26]~22_combout ),
	.A_wr_data_unfiltered_20(\A_wr_data_unfiltered[20]~23_combout ),
	.A_wr_data_unfiltered_19(\A_wr_data_unfiltered[19]~24_combout ),
	.A_wr_data_unfiltered_17(\A_wr_data_unfiltered[17]~25_combout ),
	.A_wr_data_unfiltered_30(\A_wr_data_unfiltered[30]~26_combout ),
	.A_wr_data_unfiltered_18(\A_wr_data_unfiltered[18]~27_combout ),
	.A_wr_data_unfiltered_16(\A_wr_data_unfiltered[16]~28_combout ),
	.A_wr_data_unfiltered_15(\A_wr_data_unfiltered[15]~29_combout ),
	.A_wr_data_unfiltered_12(\A_wr_data_unfiltered[12]~30_combout ),
	.A_wr_data_unfiltered_13(\A_wr_data_unfiltered[13]~31_combout ),
	.A_wr_data_unfiltered_14(\A_wr_data_unfiltered[14]~32_combout ),
	.A_wr_data_unfiltered_29(\A_wr_data_unfiltered[29]~33_combout ),
	.A_wr_dst_reg(\A_wr_dst_reg~0_combout ),
	.A_dst_regnum(\A_dst_regnum~0_combout ),
	.A_dst_regnum1(\A_dst_regnum~1_combout ),
	.A_dst_regnum2(\A_dst_regnum~2_combout ),
	.A_dst_regnum3(\A_dst_regnum~3_combout ),
	.A_dst_regnum4(\A_dst_regnum~4_combout ),
	.rf_a_rd_port_addr_0(\rf_a_rd_port_addr[0]~0_combout ),
	.rf_a_rd_port_addr_1(\rf_a_rd_port_addr[1]~1_combout ),
	.rf_a_rd_port_addr_2(\rf_a_rd_port_addr[2]~2_combout ),
	.rf_a_rd_port_addr_3(\rf_a_rd_port_addr[3]~3_combout ),
	.rf_a_rd_port_addr_4(\rf_a_rd_port_addr[4]~4_combout ),
	.clk_clk(clk_clk));

first_nios2_system_first_nios2_system_cpu_cpu_bht_module first_nios2_system_cpu_cpu_bht(
	.q_b_1(\first_nios2_system_cpu_cpu_bht|the_altsyncram|auto_generated|q_b[1] ),
	.q_b_0(\first_nios2_system_cpu_cpu_bht|the_altsyncram|auto_generated|q_b[0] ),
	.F_stall(\F_stall~0_combout ),
	.M_bht_wr_en_unfiltered(\M_bht_wr_en_unfiltered~combout ),
	.M_bht_wr_data_unfiltered_1(\M_bht_wr_data_unfiltered[1]~0_combout ),
	.M_bht_ptr_unfiltered_0(\M_bht_ptr_unfiltered[0]~q ),
	.M_bht_ptr_unfiltered_1(\M_bht_ptr_unfiltered[1]~q ),
	.M_bht_ptr_unfiltered_2(\M_bht_ptr_unfiltered[2]~q ),
	.M_bht_ptr_unfiltered_3(\M_bht_ptr_unfiltered[3]~q ),
	.M_bht_ptr_unfiltered_4(\M_bht_ptr_unfiltered[4]~q ),
	.M_bht_ptr_unfiltered_5(\M_bht_ptr_unfiltered[5]~q ),
	.M_bht_ptr_unfiltered_6(\M_bht_ptr_unfiltered[6]~q ),
	.M_bht_ptr_unfiltered_7(\M_bht_ptr_unfiltered[7]~q ),
	.F_bht_ptr_nxt_0(\F_bht_ptr_nxt[0]~combout ),
	.F_bht_ptr_nxt_1(\F_bht_ptr_nxt[1]~combout ),
	.F_bht_ptr_nxt_2(\F_bht_ptr_nxt[2]~combout ),
	.F_bht_ptr_nxt_3(\F_bht_ptr_nxt[3]~combout ),
	.F_bht_ptr_nxt_4(\F_bht_ptr_nxt[4]~combout ),
	.F_bht_ptr_nxt_5(\F_bht_ptr_nxt[5]~combout ),
	.F_bht_ptr_nxt_6(\F_bht_ptr_nxt[6]~combout ),
	.F_bht_ptr_nxt_7(\F_bht_ptr_nxt[7]~combout ),
	.M_br_mispredict(\M_br_mispredict~_wirecell_combout ),
	.clk_clk(clk_clk));

first_nios2_system_first_nios2_system_cpu_cpu_ic_tag_module first_nios2_system_cpu_cpu_ic_tag(
	.q_b_5(\first_nios2_system_cpu_cpu_ic_tag|the_altsyncram|auto_generated|q_b[5] ),
	.q_b_0(\first_nios2_system_cpu_cpu_ic_tag|the_altsyncram|auto_generated|q_b[0] ),
	.q_b_1(\first_nios2_system_cpu_cpu_ic_tag|the_altsyncram|auto_generated|q_b[1] ),
	.q_b_2(\first_nios2_system_cpu_cpu_ic_tag|the_altsyncram|auto_generated|q_b[2] ),
	.q_b_3(\first_nios2_system_cpu_cpu_ic_tag|the_altsyncram|auto_generated|q_b[3] ),
	.q_b_4(\first_nios2_system_cpu_cpu_ic_tag|the_altsyncram|auto_generated|q_b[4] ),
	.q_b_11(\first_nios2_system_cpu_cpu_ic_tag|the_altsyncram|auto_generated|q_b[11] ),
	.q_b_13(\first_nios2_system_cpu_cpu_ic_tag|the_altsyncram|auto_generated|q_b[13] ),
	.q_b_10(\first_nios2_system_cpu_cpu_ic_tag|the_altsyncram|auto_generated|q_b[10] ),
	.q_b_12(\first_nios2_system_cpu_cpu_ic_tag|the_altsyncram|auto_generated|q_b[12] ),
	.ic_tag_wraddress_0(\ic_tag_wraddress[0]~q ),
	.ic_tag_wraddress_1(\ic_tag_wraddress[1]~q ),
	.ic_tag_wraddress_2(\ic_tag_wraddress[2]~q ),
	.ic_tag_wraddress_3(\ic_tag_wraddress[3]~q ),
	.ic_tag_wraddress_4(\ic_tag_wraddress[4]~q ),
	.ic_tag_wraddress_5(\ic_tag_wraddress[5]~q ),
	.ic_fill_valid_bits_5(\ic_fill_valid_bits[5]~q ),
	.ic_fill_valid_bits_7(\ic_fill_valid_bits[7]~q ),
	.ic_fill_valid_bits_4(\ic_fill_valid_bits[4]~q ),
	.q_b_7(\first_nios2_system_cpu_cpu_ic_tag|the_altsyncram|auto_generated|q_b[7] ),
	.q_b_9(\first_nios2_system_cpu_cpu_ic_tag|the_altsyncram|auto_generated|q_b[9] ),
	.q_b_6(\first_nios2_system_cpu_cpu_ic_tag|the_altsyncram|auto_generated|q_b[6] ),
	.q_b_8(\first_nios2_system_cpu_cpu_ic_tag|the_altsyncram|auto_generated|q_b[8] ),
	.ic_fill_valid_bits_6(\ic_fill_valid_bits[6]~q ),
	.ic_fill_valid_bits_1(\ic_fill_valid_bits[1]~q ),
	.ic_fill_valid_bits_3(\ic_fill_valid_bits[3]~q ),
	.ic_fill_valid_bits_0(\ic_fill_valid_bits[0]~q ),
	.ic_fill_valid_bits_2(\ic_fill_valid_bits[2]~q ),
	.ic_fill_tag_5(ic_fill_tag_5),
	.ic_fill_tag_4(ic_fill_tag_4),
	.ic_fill_tag_3(ic_fill_tag_3),
	.ic_fill_tag_2(ic_fill_tag_2),
	.ic_fill_tag_1(ic_fill_tag_1),
	.ic_fill_tag_0(ic_fill_tag_0),
	.F_stall(\F_stall~0_combout ),
	.F_ic_tag_rd_addr_nxt_0(\F_ic_tag_rd_addr_nxt[0]~5_combout ),
	.F_ic_tag_rd_addr_nxt_1(\F_ic_tag_rd_addr_nxt[1]~7_combout ),
	.F_ic_tag_rd_addr_nxt_2(\F_ic_tag_rd_addr_nxt[2]~9_combout ),
	.F_ic_tag_rd_addr_nxt_3(\F_ic_tag_rd_addr_nxt[3]~11_combout ),
	.F_ic_tag_rd_addr_nxt_4(\F_ic_tag_rd_addr_nxt[4]~13_combout ),
	.F_ic_tag_rd_addr_nxt_5(\F_ic_tag_rd_addr_nxt[5]~15_combout ),
	.ic_tag_wren(\ic_tag_wren~combout ),
	.clk_clk(clk_clk));

first_nios2_system_first_nios2_system_cpu_cpu_ic_data_module first_nios2_system_cpu_cpu_ic_data(
	.q_b_26(\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[26] ),
	.q_b_25(\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[25] ),
	.q_b_24(\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[24] ),
	.q_b_23(\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[23] ),
	.q_b_22(\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[22] ),
	.q_b_1(\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[1] ),
	.q_b_0(\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[0] ),
	.q_b_2(\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[2] ),
	.q_b_3(\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[3] ),
	.q_b_4(\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[4] ),
	.q_b_5(\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[5] ),
	.q_b_28(\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[28] ),
	.q_b_31(\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[31] ),
	.q_b_27(\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[27] ),
	.q_b_29(\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[29] ),
	.q_b_30(\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[30] ),
	.q_b_11(\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[11] ),
	.q_b_12(\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[12] ),
	.q_b_13(\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[13] ),
	.q_b_14(\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[14] ),
	.q_b_15(\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[15] ),
	.q_b_16(\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[16] ),
	.q_b_9(\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[9] ),
	.q_b_21(\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[21] ),
	.q_b_6(\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[6] ),
	.q_b_8(\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[8] ),
	.q_b_17(\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[17] ),
	.q_b_18(\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[18] ),
	.q_b_10(\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[10] ),
	.q_b_7(\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[7] ),
	.q_b_20(\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[20] ),
	.q_b_19(\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[19] ),
	.ic_fill_line_0(ic_fill_line_0),
	.ic_fill_line_5(ic_fill_line_5),
	.ic_fill_line_4(ic_fill_line_4),
	.ic_fill_line_3(ic_fill_line_3),
	.ic_fill_line_2(ic_fill_line_2),
	.ic_fill_line_1(ic_fill_line_1),
	.F_stall(\F_stall~0_combout ),
	.ic_fill_dp_offset_0(\ic_fill_dp_offset[0]~q ),
	.ic_fill_dp_offset_1(\ic_fill_dp_offset[1]~q ),
	.ic_fill_dp_offset_2(\ic_fill_dp_offset[2]~q ),
	.i_readdatavalid_d1(\i_readdatavalid_d1~q ),
	.i_readdata_d1_26(\i_readdata_d1[26]~q ),
	.F_ic_data_rd_addr_nxt_0(\F_ic_data_rd_addr_nxt[0]~1_combout ),
	.F_ic_data_rd_addr_nxt_1(\F_ic_data_rd_addr_nxt[1]~3_combout ),
	.F_ic_data_rd_addr_nxt_2(\F_ic_data_rd_addr_nxt[2]~5_combout ),
	.F_ic_tag_rd_addr_nxt_0(\F_ic_tag_rd_addr_nxt[0]~5_combout ),
	.F_ic_tag_rd_addr_nxt_1(\F_ic_tag_rd_addr_nxt[1]~7_combout ),
	.F_ic_tag_rd_addr_nxt_2(\F_ic_tag_rd_addr_nxt[2]~9_combout ),
	.F_ic_tag_rd_addr_nxt_3(\F_ic_tag_rd_addr_nxt[3]~11_combout ),
	.F_ic_tag_rd_addr_nxt_4(\F_ic_tag_rd_addr_nxt[4]~13_combout ),
	.F_ic_tag_rd_addr_nxt_5(\F_ic_tag_rd_addr_nxt[5]~15_combout ),
	.i_readdata_d1_25(\i_readdata_d1[25]~q ),
	.i_readdata_d1_24(\i_readdata_d1[24]~q ),
	.i_readdata_d1_23(\i_readdata_d1[23]~q ),
	.i_readdata_d1_22(\i_readdata_d1[22]~q ),
	.i_readdata_d1_1(\i_readdata_d1[1]~q ),
	.i_readdata_d1_0(\i_readdata_d1[0]~q ),
	.i_readdata_d1_2(\i_readdata_d1[2]~q ),
	.i_readdata_d1_3(\i_readdata_d1[3]~q ),
	.i_readdata_d1_4(\i_readdata_d1[4]~q ),
	.i_readdata_d1_5(\i_readdata_d1[5]~q ),
	.i_readdata_d1_28(\i_readdata_d1[28]~q ),
	.i_readdata_d1_31(\i_readdata_d1[31]~q ),
	.i_readdata_d1_27(\i_readdata_d1[27]~q ),
	.i_readdata_d1_29(\i_readdata_d1[29]~q ),
	.i_readdata_d1_30(\i_readdata_d1[30]~q ),
	.i_readdata_d1_11(\i_readdata_d1[11]~q ),
	.i_readdata_d1_12(\i_readdata_d1[12]~q ),
	.i_readdata_d1_13(\i_readdata_d1[13]~q ),
	.i_readdata_d1_14(\i_readdata_d1[14]~q ),
	.i_readdata_d1_15(\i_readdata_d1[15]~q ),
	.i_readdata_d1_16(\i_readdata_d1[16]~q ),
	.i_readdata_d1_9(\i_readdata_d1[9]~q ),
	.i_readdata_d1_21(\i_readdata_d1[21]~q ),
	.i_readdata_d1_6(\i_readdata_d1[6]~q ),
	.i_readdata_d1_8(\i_readdata_d1[8]~q ),
	.i_readdata_d1_17(\i_readdata_d1[17]~q ),
	.i_readdata_d1_18(\i_readdata_d1[18]~q ),
	.i_readdata_d1_10(\i_readdata_d1[10]~q ),
	.i_readdata_d1_7(\i_readdata_d1[7]~q ),
	.i_readdata_d1_20(\i_readdata_d1[20]~q ),
	.i_readdata_d1_19(\i_readdata_d1[19]~q ),
	.clk_clk(clk_clk));

first_nios2_system_first_nios2_system_cpu_cpu_mult_cell the_first_nios2_system_cpu_cpu_mult_cell(
	.E_src1_3(\E_src1[3]~q ),
	.E_src2_22(\E_src2[22]~q ),
	.E_src1_22(\E_src1[22]~q ),
	.E_src2_23(\E_src2[23]~q ),
	.E_src1_23(\E_src1[23]~q ),
	.E_src2_24(\E_src2[24]~q ),
	.E_src1_24(\E_src1[24]~q ),
	.E_src1_0(\E_src1[0]~q ),
	.E_src2_25(\E_src2[25]~q ),
	.E_src1_25(\E_src1[25]~q ),
	.E_src1_2(\E_src1[2]~q ),
	.E_src1_31(\E_src1[31]~q ),
	.E_src2_7(\E_src2[7]~q ),
	.E_src1_7(\E_src1[7]~q ),
	.E_src2_21(\E_src2[21]~q ),
	.E_src1_21(\E_src1[21]~q ),
	.E_src2_11(\E_src2[11]~q ),
	.E_src1_11(\E_src1[11]~q ),
	.E_src2_28(\E_src2[28]~q ),
	.E_src1_28(\E_src1[28]~q ),
	.E_src2_10(\E_src2[10]~q ),
	.E_src1_10(\E_src1[10]~q ),
	.E_src2_27(\E_src2[27]~q ),
	.E_src1_27(\E_src1[27]~q ),
	.E_src2_8(\E_src2[8]~q ),
	.E_src1_8(\E_src1[8]~q ),
	.E_src2_9(\E_src2[9]~q ),
	.E_src1_9(\E_src1[9]~q ),
	.E_src1_4(\E_src1[4]~q ),
	.E_src2_5(\E_src2[5]~q ),
	.E_src1_5(\E_src1[5]~q ),
	.E_src2_6(\E_src2[6]~q ),
	.E_src1_6(\E_src1[6]~q ),
	.E_src2_26(\E_src2[26]~q ),
	.E_src1_26(\E_src1[26]~q ),
	.E_src2_20(\E_src2[20]~q ),
	.E_src1_20(\E_src1[20]~q ),
	.E_src2_19(\E_src2[19]~q ),
	.E_src1_19(\E_src1[19]~q ),
	.E_src2_17(\E_src2[17]~q ),
	.E_src1_17(\E_src1[17]~q ),
	.E_src2_30(\E_src2[30]~q ),
	.E_src1_30(\E_src1[30]~q ),
	.E_src1_1(\E_src1[1]~q ),
	.E_src2_18(\E_src2[18]~q ),
	.E_src1_18(\E_src1[18]~q ),
	.E_src2_16(\E_src2[16]~q ),
	.E_src1_16(\E_src1[16]~q ),
	.E_src2_15(\E_src2[15]~q ),
	.E_src1_15(\E_src1[15]~q ),
	.E_src2_12(\E_src2[12]~q ),
	.E_src1_12(\E_src1[12]~q ),
	.E_src2_13(\E_src2[13]~q ),
	.E_src1_13(\E_src1[13]~q ),
	.E_src2_14(\E_src2[14]~q ),
	.E_src1_14(\E_src1[14]~q ),
	.E_src2_29(\E_src2[29]~q ),
	.E_src1_29(\E_src1[29]~q ),
	.r_sync_rst(r_sync_rst),
	.A_mem_stall(\A_mem_stall~q ),
	.E_src2_3(\E_src2[3]~q ),
	.E_src2_0(\E_src2[0]~q ),
	.E_src2_2(\E_src2[2]~q ),
	.E_src2_31(\E_src2[31]~q ),
	.E_src2_4(\E_src2[4]~q ),
	.E_src2_1(\E_src2[1]~q ),
	.data_out_wire_0(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[0]~q ),
	.data_out_wire_1(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[1]~q ),
	.data_out_wire_2(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[2]~q ),
	.data_out_wire_3(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[3]~q ),
	.data_out_wire_4(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[4]~q ),
	.data_out_wire_5(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[5]~q ),
	.data_out_wire_6(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[6]~q ),
	.data_out_wire_7(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[7]~q ),
	.data_out_wire_11(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[11]~q ),
	.data_out_wire_10(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[10]~q ),
	.data_out_wire_8(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[8]~q ),
	.data_out_wire_9(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[9]~q ),
	.data_out_wire_15(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[15]~q ),
	.data_out_wire_12(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[12]~q ),
	.data_out_wire_13(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[13]~q ),
	.data_out_wire_14(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[14]~q ),
	.data_out_wire_61(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p3|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[6]~q ),
	.data_out_wire_71(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p3|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[7]~q ),
	.data_out_wire_81(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p3|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[8]~q ),
	.data_out_wire_91(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p3|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[9]~q ),
	.data_out_wire_151(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p3|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[15]~q ),
	.data_out_wire_51(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p3|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[5]~q ),
	.data_out_wire_121(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p3|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[12]~q ),
	.data_out_wire_111(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p3|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[11]~q ),
	.data_out_wire_101(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p3|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[10]~q ),
	.data_out_wire_41(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p3|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[4]~q ),
	.data_out_wire_31(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p3|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[3]~q ),
	.data_out_wire_16(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p3|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[1]~q ),
	.data_out_wire_141(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p3|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[14]~q ),
	.data_out_wire_21(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p3|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[2]~q ),
	.data_out_wire_01(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p3|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[0]~q ),
	.data_out_wire_131(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p3|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[13]~q ),
	.data_out_wire_62(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[6]~q ),
	.data_out_wire_22(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[22]~q ),
	.data_out_wire_72(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[7]~q ),
	.data_out_wire_23(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[23]~q ),
	.data_out_wire_82(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[8]~q ),
	.data_out_wire_24(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[24]~q ),
	.data_out_wire_92(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[9]~q ),
	.data_out_wire_25(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[25]~q ),
	.data_out_wire_152(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[15]~q ),
	.data_out_wire_311(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[31]~q ),
	.data_out_wire_52(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[5]~q ),
	.data_out_wire_211(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[21]~q ),
	.data_out_wire_122(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[12]~q ),
	.data_out_wire_28(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[28]~q ),
	.data_out_wire_112(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[11]~q ),
	.data_out_wire_27(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[27]~q ),
	.data_out_wire_102(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[10]~q ),
	.data_out_wire_26(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[26]~q ),
	.data_out_wire_42(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[4]~q ),
	.data_out_wire_20(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[20]~q ),
	.data_out_wire_32(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[3]~q ),
	.data_out_wire_19(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[19]~q ),
	.data_out_wire_17(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[1]~q ),
	.data_out_wire_171(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[17]~q ),
	.data_out_wire_142(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[14]~q ),
	.data_out_wire_30(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[30]~q ),
	.data_out_wire_29(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[2]~q ),
	.data_out_wire_18(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[18]~q ),
	.data_out_wire_02(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[0]~q ),
	.data_out_wire_161(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[16]~q ),
	.data_out_wire_132(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[13]~q ),
	.data_out_wire_291(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[29]~q ),
	.clk_clk(clk_clk));

first_nios2_system_first_nios2_system_cpu_cpu_register_bank_b_module first_nios2_system_cpu_cpu_register_bank_b(
	.q_b_0(\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[0] ),
	.q_b_1(\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[1] ),
	.q_b_2(\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[2] ),
	.q_b_3(\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[3] ),
	.q_b_4(\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[4] ),
	.q_b_5(\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[5] ),
	.q_b_6(\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[6] ),
	.q_b_7(\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[7] ),
	.q_b_22(\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[22] ),
	.q_b_23(\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[23] ),
	.q_b_24(\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[24] ),
	.q_b_25(\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[25] ),
	.q_b_31(\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[31] ),
	.q_b_21(\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[21] ),
	.q_b_11(\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[11] ),
	.q_b_28(\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[28] ),
	.q_b_10(\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[10] ),
	.q_b_27(\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[27] ),
	.q_b_8(\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[8] ),
	.q_b_9(\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[9] ),
	.q_b_26(\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[26] ),
	.q_b_20(\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[20] ),
	.q_b_19(\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[19] ),
	.q_b_17(\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[17] ),
	.q_b_30(\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[30] ),
	.q_b_18(\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[18] ),
	.q_b_16(\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[16] ),
	.q_b_15(\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[15] ),
	.q_b_12(\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[12] ),
	.q_b_13(\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[13] ),
	.q_b_14(\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[14] ),
	.q_b_29(\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[29] ),
	.A_wr_data_unfiltered_0(\A_wr_data_unfiltered[0]~2_combout ),
	.A_wr_data_unfiltered_1(\A_wr_data_unfiltered[1]~3_combout ),
	.A_wr_data_unfiltered_2(\A_wr_data_unfiltered[2]~4_combout ),
	.A_wr_data_unfiltered_3(\A_wr_data_unfiltered[3]~5_combout ),
	.A_wr_data_unfiltered_4(\A_wr_data_unfiltered[4]~6_combout ),
	.A_wr_data_unfiltered_5(\A_wr_data_unfiltered[5]~7_combout ),
	.A_wr_data_unfiltered_6(\A_wr_data_unfiltered[6]~8_combout ),
	.A_wr_data_unfiltered_7(\A_wr_data_unfiltered[7]~9_combout ),
	.A_wr_data_unfiltered_22(\A_wr_data_unfiltered[22]~10_combout ),
	.A_wr_data_unfiltered_23(\A_wr_data_unfiltered[23]~11_combout ),
	.A_wr_data_unfiltered_24(\A_wr_data_unfiltered[24]~12_combout ),
	.A_wr_data_unfiltered_25(\A_wr_data_unfiltered[25]~13_combout ),
	.A_wr_data_unfiltered_31(\A_wr_data_unfiltered[31]~14_combout ),
	.A_wr_data_unfiltered_21(\A_wr_data_unfiltered[21]~15_combout ),
	.A_wr_data_unfiltered_11(\A_wr_data_unfiltered[11]~16_combout ),
	.A_wr_data_unfiltered_28(\A_wr_data_unfiltered[28]~17_combout ),
	.A_wr_data_unfiltered_10(\A_wr_data_unfiltered[10]~18_combout ),
	.A_wr_data_unfiltered_27(\A_wr_data_unfiltered[27]~19_combout ),
	.A_wr_data_unfiltered_8(\A_wr_data_unfiltered[8]~20_combout ),
	.A_wr_data_unfiltered_9(\A_wr_data_unfiltered[9]~21_combout ),
	.A_wr_data_unfiltered_26(\A_wr_data_unfiltered[26]~22_combout ),
	.A_wr_data_unfiltered_20(\A_wr_data_unfiltered[20]~23_combout ),
	.A_wr_data_unfiltered_19(\A_wr_data_unfiltered[19]~24_combout ),
	.A_wr_data_unfiltered_17(\A_wr_data_unfiltered[17]~25_combout ),
	.A_wr_data_unfiltered_30(\A_wr_data_unfiltered[30]~26_combout ),
	.A_wr_data_unfiltered_18(\A_wr_data_unfiltered[18]~27_combout ),
	.A_wr_data_unfiltered_16(\A_wr_data_unfiltered[16]~28_combout ),
	.A_wr_data_unfiltered_15(\A_wr_data_unfiltered[15]~29_combout ),
	.A_wr_data_unfiltered_12(\A_wr_data_unfiltered[12]~30_combout ),
	.A_wr_data_unfiltered_13(\A_wr_data_unfiltered[13]~31_combout ),
	.A_wr_data_unfiltered_14(\A_wr_data_unfiltered[14]~32_combout ),
	.A_wr_data_unfiltered_29(\A_wr_data_unfiltered[29]~33_combout ),
	.A_wr_dst_reg(\A_wr_dst_reg~0_combout ),
	.A_dst_regnum(\A_dst_regnum~0_combout ),
	.A_dst_regnum1(\A_dst_regnum~1_combout ),
	.A_dst_regnum2(\A_dst_regnum~2_combout ),
	.A_dst_regnum3(\A_dst_regnum~3_combout ),
	.A_dst_regnum4(\A_dst_regnum~4_combout ),
	.rf_b_rd_port_addr_0(\rf_b_rd_port_addr[0]~0_combout ),
	.rf_b_rd_port_addr_1(\rf_b_rd_port_addr[1]~1_combout ),
	.rf_b_rd_port_addr_2(\rf_b_rd_port_addr[2]~2_combout ),
	.rf_b_rd_port_addr_3(\rf_b_rd_port_addr[3]~3_combout ),
	.rf_b_rd_port_addr_4(\rf_b_rd_port_addr[4]~4_combout ),
	.clk_clk(clk_clk));

first_nios2_system_first_nios2_system_cpu_cpu_nios2_oci the_first_nios2_system_cpu_cpu_nios2_oci(
	.readdata_0(readdata_0),
	.readdata_1(readdata_1),
	.readdata_2(readdata_2),
	.readdata_3(readdata_3),
	.readdata_4(readdata_4),
	.readdata_5(readdata_5),
	.readdata_6(readdata_6),
	.readdata_7(readdata_7),
	.readdata_22(readdata_22),
	.readdata_23(readdata_23),
	.readdata_24(readdata_24),
	.readdata_25(readdata_25),
	.readdata_31(readdata_31),
	.readdata_21(readdata_21),
	.readdata_11(readdata_11),
	.readdata_28(readdata_28),
	.readdata_10(readdata_10),
	.readdata_27(readdata_27),
	.readdata_8(readdata_8),
	.readdata_9(readdata_9),
	.readdata_26(readdata_26),
	.readdata_20(readdata_20),
	.readdata_19(readdata_19),
	.readdata_17(readdata_17),
	.readdata_30(readdata_30),
	.readdata_18(readdata_18),
	.readdata_16(readdata_16),
	.readdata_15(readdata_15),
	.readdata_12(readdata_12),
	.readdata_13(readdata_13),
	.readdata_14(readdata_14),
	.readdata_29(readdata_29),
	.sr_0(sr_0),
	.ir_out_0(ir_out_0),
	.ir_out_1(ir_out_1),
	.d_write(d_write1),
	.r_sync_rst(r_sync_rst),
	.W_debug_mode(W_debug_mode1),
	.oci_single_step_mode(\the_first_nios2_system_cpu_cpu_nios2_oci|the_first_nios2_system_cpu_cpu_nios2_avalon_reg|oci_single_step_mode~q ),
	.jtag_break(\the_first_nios2_system_cpu_cpu_nios2_oci|the_first_nios2_system_cpu_cpu_nios2_oci_debug|jtag_break~q ),
	.saved_grant_0(saved_grant_0),
	.waitrequest(debug_mem_slave_waitrequest),
	.mem_used_1(mem_used_1),
	.WideOr1(WideOr14),
	.mem(mem),
	.oci_ienable_1(\the_first_nios2_system_cpu_cpu_nios2_oci|the_first_nios2_system_cpu_cpu_nios2_avalon_reg|oci_ienable[1]~q ),
	.oci_ienable_16(\the_first_nios2_system_cpu_cpu_nios2_oci|the_first_nios2_system_cpu_cpu_nios2_avalon_reg|oci_ienable[16]~q ),
	.writedata_nxt({src_payload34,src_payload40,src_payload45,src_payload36,src_payload31,src_payload30,src_payload29,src_payload28,src_payload33,src_payload32,src_payload21,src_payload19,src_payload20,src_payload22,src_payload23,src_payload17,src_payload41,src_payload44,src_payload43,
src_payload42,src_payload35,src_payload37,src_payload39,src_payload38,src_payload27,src_payload26,src_payload25,src_payload24,src_payload,src_payload18,src_payload16,src_payload3}),
	.address_nxt({src_data_46,src_data_45,src_data_44,src_data_43,src_data_42,src_data_41,src_data_40,src_data_39,src_data_38}),
	.debugaccess_nxt(src_payload1),
	.r_early_rst(r_early_rst),
	.byteenable_nxt({src_data_35,src_data_34,src_data_33,src_data_32}),
	.altera_internal_jtag(altera_internal_jtag),
	.altera_internal_jtag1(altera_internal_jtag1),
	.state_1(state_1),
	.state_4(state_4),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.state_8(state_8),
	.splitter_nodes_receive_1_3(splitter_nodes_receive_1_3),
	.irf_reg_0_2(irf_reg_0_2),
	.irf_reg_1_2(irf_reg_1_2),
	.clk_clk(clk_clk));

dffeas \ic_tag_wraddress[0] (
	.clk(clk_clk),
	.d(\ic_tag_wraddress_nxt~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(!clr_break_line1),
	.ena(vcc),
	.q(\ic_tag_wraddress[0]~q ),
	.prn(vcc));
defparam \ic_tag_wraddress[0] .is_wysiwyg = "true";
defparam \ic_tag_wraddress[0] .power_up = "low";

dffeas \ic_tag_wraddress[1] (
	.clk(clk_clk),
	.d(\ic_tag_wraddress_nxt[1]~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(!clr_break_line1),
	.sload(gnd),
	.ena(vcc),
	.q(\ic_tag_wraddress[1]~q ),
	.prn(vcc));
defparam \ic_tag_wraddress[1] .is_wysiwyg = "true";
defparam \ic_tag_wraddress[1] .power_up = "low";

dffeas \ic_tag_wraddress[2] (
	.clk(clk_clk),
	.d(\ic_tag_wraddress_nxt[2]~8_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(!clr_break_line1),
	.sload(gnd),
	.ena(vcc),
	.q(\ic_tag_wraddress[2]~q ),
	.prn(vcc));
defparam \ic_tag_wraddress[2] .is_wysiwyg = "true";
defparam \ic_tag_wraddress[2] .power_up = "low";

dffeas \ic_tag_wraddress[3] (
	.clk(clk_clk),
	.d(\ic_tag_wraddress_nxt[3]~9_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(!clr_break_line1),
	.sload(gnd),
	.ena(vcc),
	.q(\ic_tag_wraddress[3]~q ),
	.prn(vcc));
defparam \ic_tag_wraddress[3] .is_wysiwyg = "true";
defparam \ic_tag_wraddress[3] .power_up = "low";

dffeas \ic_tag_wraddress[4] (
	.clk(clk_clk),
	.d(\ic_tag_wraddress_nxt[4]~10_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(!clr_break_line1),
	.sload(gnd),
	.ena(vcc),
	.q(\ic_tag_wraddress[4]~q ),
	.prn(vcc));
defparam \ic_tag_wraddress[4] .is_wysiwyg = "true";
defparam \ic_tag_wraddress[4] .power_up = "low";

dffeas \ic_tag_wraddress[5] (
	.clk(clk_clk),
	.d(\ic_tag_wraddress_nxt[5]~11_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(!clr_break_line1),
	.sload(gnd),
	.ena(vcc),
	.q(\ic_tag_wraddress[5]~q ),
	.prn(vcc));
defparam \ic_tag_wraddress[5] .is_wysiwyg = "true";
defparam \ic_tag_wraddress[5] .power_up = "low";

dffeas \ic_fill_valid_bits[5] (
	.clk(clk_clk),
	.d(\ic_fill_valid_bits_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\ic_tag_clr_valid_bits_nxt~combout ),
	.sload(gnd),
	.ena(\ic_fill_valid_bits_en~combout ),
	.q(\ic_fill_valid_bits[5]~q ),
	.prn(vcc));
defparam \ic_fill_valid_bits[5] .is_wysiwyg = "true";
defparam \ic_fill_valid_bits[5] .power_up = "low";

dffeas \ic_fill_valid_bits[7] (
	.clk(clk_clk),
	.d(\ic_fill_valid_bits_nxt~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\ic_tag_clr_valid_bits_nxt~combout ),
	.sload(gnd),
	.ena(\ic_fill_valid_bits_en~combout ),
	.q(\ic_fill_valid_bits[7]~q ),
	.prn(vcc));
defparam \ic_fill_valid_bits[7] .is_wysiwyg = "true";
defparam \ic_fill_valid_bits[7] .power_up = "low";

dffeas \ic_fill_valid_bits[4] (
	.clk(clk_clk),
	.d(\ic_fill_valid_bits_nxt~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\ic_tag_clr_valid_bits_nxt~combout ),
	.sload(gnd),
	.ena(\ic_fill_valid_bits_en~combout ),
	.q(\ic_fill_valid_bits[4]~q ),
	.prn(vcc));
defparam \ic_fill_valid_bits[4] .is_wysiwyg = "true";
defparam \ic_fill_valid_bits[4] .power_up = "low";

dffeas \ic_fill_valid_bits[6] (
	.clk(clk_clk),
	.d(\ic_fill_valid_bits_nxt~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\ic_tag_clr_valid_bits_nxt~combout ),
	.sload(gnd),
	.ena(\ic_fill_valid_bits_en~combout ),
	.q(\ic_fill_valid_bits[6]~q ),
	.prn(vcc));
defparam \ic_fill_valid_bits[6] .is_wysiwyg = "true";
defparam \ic_fill_valid_bits[6] .power_up = "low";

dffeas \ic_fill_valid_bits[1] (
	.clk(clk_clk),
	.d(\ic_fill_valid_bits_nxt~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\ic_tag_clr_valid_bits_nxt~combout ),
	.sload(gnd),
	.ena(\ic_fill_valid_bits_en~combout ),
	.q(\ic_fill_valid_bits[1]~q ),
	.prn(vcc));
defparam \ic_fill_valid_bits[1] .is_wysiwyg = "true";
defparam \ic_fill_valid_bits[1] .power_up = "low";

dffeas \ic_fill_valid_bits[3] (
	.clk(clk_clk),
	.d(\ic_fill_valid_bits_nxt~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\ic_tag_clr_valid_bits_nxt~combout ),
	.sload(gnd),
	.ena(\ic_fill_valid_bits_en~combout ),
	.q(\ic_fill_valid_bits[3]~q ),
	.prn(vcc));
defparam \ic_fill_valid_bits[3] .is_wysiwyg = "true";
defparam \ic_fill_valid_bits[3] .power_up = "low";

dffeas \ic_fill_valid_bits[0] (
	.clk(clk_clk),
	.d(\ic_fill_valid_bits_nxt~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\ic_tag_clr_valid_bits_nxt~combout ),
	.sload(gnd),
	.ena(\ic_fill_valid_bits_en~combout ),
	.q(\ic_fill_valid_bits[0]~q ),
	.prn(vcc));
defparam \ic_fill_valid_bits[0] .is_wysiwyg = "true";
defparam \ic_fill_valid_bits[0] .power_up = "low";

dffeas \ic_fill_valid_bits[2] (
	.clk(clk_clk),
	.d(\ic_fill_valid_bits_nxt~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\ic_tag_clr_valid_bits_nxt~combout ),
	.sload(gnd),
	.ena(\ic_fill_valid_bits_en~combout ),
	.q(\ic_fill_valid_bits[2]~q ),
	.prn(vcc));
defparam \ic_fill_valid_bits[2] .is_wysiwyg = "true";
defparam \ic_fill_valid_bits[2] .power_up = "low";

cyclonev_lcell_comb \rf_b_rd_port_addr[0]~0 (
	.dataa(!\D_iw[22]~q ),
	.datab(!\F_stall~0_combout ),
	.datac(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[22] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rf_b_rd_port_addr[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rf_b_rd_port_addr[0]~0 .extended_lut = "off";
defparam \rf_b_rd_port_addr[0]~0 .lut_mask = 64'h4747474747474747;
defparam \rf_b_rd_port_addr[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \rf_b_rd_port_addr[1]~1 (
	.dataa(!\D_iw[23]~q ),
	.datab(!\F_stall~0_combout ),
	.datac(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[23] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rf_b_rd_port_addr[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rf_b_rd_port_addr[1]~1 .extended_lut = "off";
defparam \rf_b_rd_port_addr[1]~1 .lut_mask = 64'h4747474747474747;
defparam \rf_b_rd_port_addr[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \rf_b_rd_port_addr[2]~2 (
	.dataa(!\D_iw[24]~q ),
	.datab(!\F_stall~0_combout ),
	.datac(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[24] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rf_b_rd_port_addr[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rf_b_rd_port_addr[2]~2 .extended_lut = "off";
defparam \rf_b_rd_port_addr[2]~2 .lut_mask = 64'h4747474747474747;
defparam \rf_b_rd_port_addr[2]~2 .shared_arith = "off";

cyclonev_lcell_comb \rf_b_rd_port_addr[3]~3 (
	.dataa(!\D_iw[25]~q ),
	.datab(!\F_stall~0_combout ),
	.datac(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[25] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rf_b_rd_port_addr[3]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rf_b_rd_port_addr[3]~3 .extended_lut = "off";
defparam \rf_b_rd_port_addr[3]~3 .lut_mask = 64'h4747474747474747;
defparam \rf_b_rd_port_addr[3]~3 .shared_arith = "off";

cyclonev_lcell_comb \rf_b_rd_port_addr[4]~4 (
	.dataa(!\D_iw[26]~q ),
	.datab(!\F_stall~0_combout ),
	.datac(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[26] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rf_b_rd_port_addr[4]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rf_b_rd_port_addr[4]~4 .extended_lut = "off";
defparam \rf_b_rd_port_addr[4]~4 .lut_mask = 64'h4747474747474747;
defparam \rf_b_rd_port_addr[4]~4 .shared_arith = "off";

cyclonev_lcell_comb \rf_a_rd_port_addr[0]~0 (
	.dataa(!\D_iw[27]~q ),
	.datab(!\F_stall~0_combout ),
	.datac(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[27] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rf_a_rd_port_addr[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rf_a_rd_port_addr[0]~0 .extended_lut = "off";
defparam \rf_a_rd_port_addr[0]~0 .lut_mask = 64'h4747474747474747;
defparam \rf_a_rd_port_addr[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \rf_a_rd_port_addr[1]~1 (
	.dataa(!\D_iw[28]~q ),
	.datab(!\F_stall~0_combout ),
	.datac(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[28] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rf_a_rd_port_addr[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rf_a_rd_port_addr[1]~1 .extended_lut = "off";
defparam \rf_a_rd_port_addr[1]~1 .lut_mask = 64'h4747474747474747;
defparam \rf_a_rd_port_addr[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \rf_a_rd_port_addr[2]~2 (
	.dataa(!\D_iw[29]~q ),
	.datab(!\F_stall~0_combout ),
	.datac(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[29] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rf_a_rd_port_addr[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rf_a_rd_port_addr[2]~2 .extended_lut = "off";
defparam \rf_a_rd_port_addr[2]~2 .lut_mask = 64'h4747474747474747;
defparam \rf_a_rd_port_addr[2]~2 .shared_arith = "off";

cyclonev_lcell_comb \rf_a_rd_port_addr[3]~3 (
	.dataa(!\D_iw[30]~q ),
	.datab(!\F_stall~0_combout ),
	.datac(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[30] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rf_a_rd_port_addr[3]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rf_a_rd_port_addr[3]~3 .extended_lut = "off";
defparam \rf_a_rd_port_addr[3]~3 .lut_mask = 64'h4747474747474747;
defparam \rf_a_rd_port_addr[3]~3 .shared_arith = "off";

cyclonev_lcell_comb \rf_a_rd_port_addr[4]~4 (
	.dataa(!\D_iw[31]~q ),
	.datab(!\F_stall~0_combout ),
	.datac(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[31] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rf_a_rd_port_addr[4]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rf_a_rd_port_addr[4]~4 .extended_lut = "off";
defparam \rf_a_rd_port_addr[4]~4 .lut_mask = 64'h4747474747474747;
defparam \rf_a_rd_port_addr[4]~4 .shared_arith = "off";

dffeas \i_readdata_d1[26] (
	.clk(clk_clk),
	.d(i_readdata[26]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[26]~q ),
	.prn(vcc));
defparam \i_readdata_d1[26] .is_wysiwyg = "true";
defparam \i_readdata_d1[26] .power_up = "low";

dffeas \i_readdata_d1[25] (
	.clk(clk_clk),
	.d(i_readdata[25]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[25]~q ),
	.prn(vcc));
defparam \i_readdata_d1[25] .is_wysiwyg = "true";
defparam \i_readdata_d1[25] .power_up = "low";

dffeas \i_readdata_d1[24] (
	.clk(clk_clk),
	.d(i_readdata[24]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[24]~q ),
	.prn(vcc));
defparam \i_readdata_d1[24] .is_wysiwyg = "true";
defparam \i_readdata_d1[24] .power_up = "low";

dffeas \i_readdata_d1[23] (
	.clk(clk_clk),
	.d(i_readdata[23]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[23]~q ),
	.prn(vcc));
defparam \i_readdata_d1[23] .is_wysiwyg = "true";
defparam \i_readdata_d1[23] .power_up = "low";

dffeas \i_readdata_d1[22] (
	.clk(clk_clk),
	.d(i_readdata[22]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[22]~q ),
	.prn(vcc));
defparam \i_readdata_d1[22] .is_wysiwyg = "true";
defparam \i_readdata_d1[22] .power_up = "low";

dffeas \i_readdata_d1[1] (
	.clk(clk_clk),
	.d(i_readdata[1]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[1]~q ),
	.prn(vcc));
defparam \i_readdata_d1[1] .is_wysiwyg = "true";
defparam \i_readdata_d1[1] .power_up = "low";

dffeas \i_readdata_d1[0] (
	.clk(clk_clk),
	.d(i_readdata[0]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[0]~q ),
	.prn(vcc));
defparam \i_readdata_d1[0] .is_wysiwyg = "true";
defparam \i_readdata_d1[0] .power_up = "low";

dffeas \i_readdata_d1[2] (
	.clk(clk_clk),
	.d(i_readdata[2]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[2]~q ),
	.prn(vcc));
defparam \i_readdata_d1[2] .is_wysiwyg = "true";
defparam \i_readdata_d1[2] .power_up = "low";

dffeas ic_tag_clr_valid_bits(
	.clk(clk_clk),
	.d(\ic_tag_clr_valid_bits~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ic_tag_clr_valid_bits~q ),
	.prn(vcc));
defparam ic_tag_clr_valid_bits.is_wysiwyg = "true";
defparam ic_tag_clr_valid_bits.power_up = "low";

cyclonev_lcell_comb ic_tag_wren(
	.dataa(!\i_readdatavalid_d1~q ),
	.datab(!\ic_tag_clr_valid_bits~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_tag_wren~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam ic_tag_wren.extended_lut = "off";
defparam ic_tag_wren.lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam ic_tag_wren.shared_arith = "off";

dffeas \i_readdata_d1[3] (
	.clk(clk_clk),
	.d(i_readdata[3]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[3]~q ),
	.prn(vcc));
defparam \i_readdata_d1[3] .is_wysiwyg = "true";
defparam \i_readdata_d1[3] .power_up = "low";

dffeas \i_readdata_d1[4] (
	.clk(clk_clk),
	.d(i_readdata[4]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[4]~q ),
	.prn(vcc));
defparam \i_readdata_d1[4] .is_wysiwyg = "true";
defparam \i_readdata_d1[4] .power_up = "low";

dffeas \i_readdata_d1[5] (
	.clk(clk_clk),
	.d(i_readdata[5]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[5]~q ),
	.prn(vcc));
defparam \i_readdata_d1[5] .is_wysiwyg = "true";
defparam \i_readdata_d1[5] .power_up = "low";

dffeas \i_readdata_d1[28] (
	.clk(clk_clk),
	.d(i_readdata[28]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[28]~q ),
	.prn(vcc));
defparam \i_readdata_d1[28] .is_wysiwyg = "true";
defparam \i_readdata_d1[28] .power_up = "low";

dffeas \i_readdata_d1[31] (
	.clk(clk_clk),
	.d(i_readdata[31]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[31]~q ),
	.prn(vcc));
defparam \i_readdata_d1[31] .is_wysiwyg = "true";
defparam \i_readdata_d1[31] .power_up = "low";

dffeas \i_readdata_d1[27] (
	.clk(clk_clk),
	.d(i_readdata[27]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[27]~q ),
	.prn(vcc));
defparam \i_readdata_d1[27] .is_wysiwyg = "true";
defparam \i_readdata_d1[27] .power_up = "low";

dffeas \i_readdata_d1[29] (
	.clk(clk_clk),
	.d(i_readdata[29]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[29]~q ),
	.prn(vcc));
defparam \i_readdata_d1[29] .is_wysiwyg = "true";
defparam \i_readdata_d1[29] .power_up = "low";

dffeas \i_readdata_d1[30] (
	.clk(clk_clk),
	.d(i_readdata[30]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[30]~q ),
	.prn(vcc));
defparam \i_readdata_d1[30] .is_wysiwyg = "true";
defparam \i_readdata_d1[30] .power_up = "low";

dffeas \i_readdata_d1[11] (
	.clk(clk_clk),
	.d(i_readdata[11]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[11]~q ),
	.prn(vcc));
defparam \i_readdata_d1[11] .is_wysiwyg = "true";
defparam \i_readdata_d1[11] .power_up = "low";

dffeas \i_readdata_d1[12] (
	.clk(clk_clk),
	.d(i_readdata[12]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[12]~q ),
	.prn(vcc));
defparam \i_readdata_d1[12] .is_wysiwyg = "true";
defparam \i_readdata_d1[12] .power_up = "low";

dffeas \i_readdata_d1[13] (
	.clk(clk_clk),
	.d(i_readdata[13]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[13]~q ),
	.prn(vcc));
defparam \i_readdata_d1[13] .is_wysiwyg = "true";
defparam \i_readdata_d1[13] .power_up = "low";

dffeas \i_readdata_d1[14] (
	.clk(clk_clk),
	.d(i_readdata[14]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[14]~q ),
	.prn(vcc));
defparam \i_readdata_d1[14] .is_wysiwyg = "true";
defparam \i_readdata_d1[14] .power_up = "low";

dffeas \i_readdata_d1[15] (
	.clk(clk_clk),
	.d(i_readdata[15]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[15]~q ),
	.prn(vcc));
defparam \i_readdata_d1[15] .is_wysiwyg = "true";
defparam \i_readdata_d1[15] .power_up = "low";

dffeas \i_readdata_d1[16] (
	.clk(clk_clk),
	.d(i_readdata[16]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[16]~q ),
	.prn(vcc));
defparam \i_readdata_d1[16] .is_wysiwyg = "true";
defparam \i_readdata_d1[16] .power_up = "low";

dffeas \i_readdata_d1[9] (
	.clk(clk_clk),
	.d(i_readdata[9]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[9]~q ),
	.prn(vcc));
defparam \i_readdata_d1[9] .is_wysiwyg = "true";
defparam \i_readdata_d1[9] .power_up = "low";

dffeas \i_readdata_d1[21] (
	.clk(clk_clk),
	.d(i_readdata[21]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[21]~q ),
	.prn(vcc));
defparam \i_readdata_d1[21] .is_wysiwyg = "true";
defparam \i_readdata_d1[21] .power_up = "low";

dffeas \i_readdata_d1[6] (
	.clk(clk_clk),
	.d(i_readdata[6]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[6]~q ),
	.prn(vcc));
defparam \i_readdata_d1[6] .is_wysiwyg = "true";
defparam \i_readdata_d1[6] .power_up = "low";

dffeas \i_readdata_d1[8] (
	.clk(clk_clk),
	.d(i_readdata[8]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[8]~q ),
	.prn(vcc));
defparam \i_readdata_d1[8] .is_wysiwyg = "true";
defparam \i_readdata_d1[8] .power_up = "low";

dffeas \i_readdata_d1[17] (
	.clk(clk_clk),
	.d(i_readdata[17]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[17]~q ),
	.prn(vcc));
defparam \i_readdata_d1[17] .is_wysiwyg = "true";
defparam \i_readdata_d1[17] .power_up = "low";

dffeas \i_readdata_d1[18] (
	.clk(clk_clk),
	.d(i_readdata[18]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[18]~q ),
	.prn(vcc));
defparam \i_readdata_d1[18] .is_wysiwyg = "true";
defparam \i_readdata_d1[18] .power_up = "low";

dffeas \i_readdata_d1[10] (
	.clk(clk_clk),
	.d(i_readdata[10]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[10]~q ),
	.prn(vcc));
defparam \i_readdata_d1[10] .is_wysiwyg = "true";
defparam \i_readdata_d1[10] .power_up = "low";

dffeas \i_readdata_d1[7] (
	.clk(clk_clk),
	.d(i_readdata[7]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[7]~q ),
	.prn(vcc));
defparam \i_readdata_d1[7] .is_wysiwyg = "true";
defparam \i_readdata_d1[7] .power_up = "low";

dffeas \i_readdata_d1[20] (
	.clk(clk_clk),
	.d(i_readdata[20]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[20]~q ),
	.prn(vcc));
defparam \i_readdata_d1[20] .is_wysiwyg = "true";
defparam \i_readdata_d1[20] .power_up = "low";

dffeas \i_readdata_d1[19] (
	.clk(clk_clk),
	.d(i_readdata[19]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[19]~q ),
	.prn(vcc));
defparam \i_readdata_d1[19] .is_wysiwyg = "true";
defparam \i_readdata_d1[19] .power_up = "low";

dffeas M_ctrl_br_cond(
	.clk(clk_clk),
	.d(\E_ctrl_br_cond~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_ctrl_br_cond~q ),
	.prn(vcc));
defparam M_ctrl_br_cond.is_wysiwyg = "true";
defparam M_ctrl_br_cond.power_up = "low";

cyclonev_lcell_comb M_bht_wr_en_unfiltered(
	.dataa(!\M_valid_from_E~q ),
	.datab(!\M_ctrl_br_cond~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_bht_wr_en_unfiltered~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam M_bht_wr_en_unfiltered.extended_lut = "off";
defparam M_bht_wr_en_unfiltered.lut_mask = 64'h7777777777777777;
defparam M_bht_wr_en_unfiltered.shared_arith = "off";

dffeas \M_bht_data[1] (
	.clk(clk_clk),
	.d(\E_bht_data[1]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_bht_data[1]~q ),
	.prn(vcc));
defparam \M_bht_data[1] .is_wysiwyg = "true";
defparam \M_bht_data[1] .power_up = "low";

dffeas \M_bht_data[0] (
	.clk(clk_clk),
	.d(\E_bht_data[0]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_bht_data[0]~q ),
	.prn(vcc));
defparam \M_bht_data[0] .is_wysiwyg = "true";
defparam \M_bht_data[0] .power_up = "low";

dffeas M_br_mispredict(
	.clk(clk_clk),
	.d(\E_br_mispredict~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_br_mispredict~q ),
	.prn(vcc));
defparam M_br_mispredict.is_wysiwyg = "true";
defparam M_br_mispredict.power_up = "low";

cyclonev_lcell_comb \M_bht_wr_data_unfiltered[1]~0 (
	.dataa(!\M_bht_data[1]~q ),
	.datab(!\M_bht_data[0]~q ),
	.datac(!\M_br_mispredict~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_bht_wr_data_unfiltered[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_bht_wr_data_unfiltered[1]~0 .extended_lut = "off";
defparam \M_bht_wr_data_unfiltered[1]~0 .lut_mask = 64'h9696969696969696;
defparam \M_bht_wr_data_unfiltered[1]~0 .shared_arith = "off";

dffeas \M_bht_ptr_unfiltered[0] (
	.clk(clk_clk),
	.d(\E_bht_ptr[0]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_bht_ptr_unfiltered[0]~q ),
	.prn(vcc));
defparam \M_bht_ptr_unfiltered[0] .is_wysiwyg = "true";
defparam \M_bht_ptr_unfiltered[0] .power_up = "low";

dffeas \M_bht_ptr_unfiltered[1] (
	.clk(clk_clk),
	.d(\E_bht_ptr[1]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_bht_ptr_unfiltered[1]~q ),
	.prn(vcc));
defparam \M_bht_ptr_unfiltered[1] .is_wysiwyg = "true";
defparam \M_bht_ptr_unfiltered[1] .power_up = "low";

dffeas \M_bht_ptr_unfiltered[2] (
	.clk(clk_clk),
	.d(\E_bht_ptr[2]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_bht_ptr_unfiltered[2]~q ),
	.prn(vcc));
defparam \M_bht_ptr_unfiltered[2] .is_wysiwyg = "true";
defparam \M_bht_ptr_unfiltered[2] .power_up = "low";

dffeas \M_bht_ptr_unfiltered[3] (
	.clk(clk_clk),
	.d(\E_bht_ptr[3]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_bht_ptr_unfiltered[3]~q ),
	.prn(vcc));
defparam \M_bht_ptr_unfiltered[3] .is_wysiwyg = "true";
defparam \M_bht_ptr_unfiltered[3] .power_up = "low";

dffeas \M_bht_ptr_unfiltered[4] (
	.clk(clk_clk),
	.d(\E_bht_ptr[4]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_bht_ptr_unfiltered[4]~q ),
	.prn(vcc));
defparam \M_bht_ptr_unfiltered[4] .is_wysiwyg = "true";
defparam \M_bht_ptr_unfiltered[4] .power_up = "low";

dffeas \M_bht_ptr_unfiltered[5] (
	.clk(clk_clk),
	.d(\E_bht_ptr[5]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_bht_ptr_unfiltered[5]~q ),
	.prn(vcc));
defparam \M_bht_ptr_unfiltered[5] .is_wysiwyg = "true";
defparam \M_bht_ptr_unfiltered[5] .power_up = "low";

dffeas \M_bht_ptr_unfiltered[6] (
	.clk(clk_clk),
	.d(\E_bht_ptr[6]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_bht_ptr_unfiltered[6]~q ),
	.prn(vcc));
defparam \M_bht_ptr_unfiltered[6] .is_wysiwyg = "true";
defparam \M_bht_ptr_unfiltered[6] .power_up = "low";

dffeas \M_bht_ptr_unfiltered[7] (
	.clk(clk_clk),
	.d(\E_bht_ptr[7]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_bht_ptr_unfiltered[7]~q ),
	.prn(vcc));
defparam \M_bht_ptr_unfiltered[7] .is_wysiwyg = "true";
defparam \M_bht_ptr_unfiltered[7] .power_up = "low";

dffeas \M_br_cond_taken_history[0] (
	.clk(clk_clk),
	.d(\E_br_result~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\M_br_cond_taken_history[0]~0_combout ),
	.q(\M_br_cond_taken_history[0]~q ),
	.prn(vcc));
defparam \M_br_cond_taken_history[0] .is_wysiwyg = "true";
defparam \M_br_cond_taken_history[0] .power_up = "low";

cyclonev_lcell_comb \F_bht_ptr_nxt[0] (
	.dataa(!\F_ic_data_rd_addr_nxt[0]~1_combout ),
	.datab(!\M_br_cond_taken_history[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_bht_ptr_nxt[0]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_bht_ptr_nxt[0] .extended_lut = "off";
defparam \F_bht_ptr_nxt[0] .lut_mask = 64'h6666666666666666;
defparam \F_bht_ptr_nxt[0] .shared_arith = "off";

dffeas \M_br_cond_taken_history[1] (
	.clk(clk_clk),
	.d(\M_br_cond_taken_history[0]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\M_br_cond_taken_history[0]~0_combout ),
	.q(\M_br_cond_taken_history[1]~q ),
	.prn(vcc));
defparam \M_br_cond_taken_history[1] .is_wysiwyg = "true";
defparam \M_br_cond_taken_history[1] .power_up = "low";

cyclonev_lcell_comb \F_bht_ptr_nxt[1] (
	.dataa(!\F_ic_data_rd_addr_nxt[1]~3_combout ),
	.datab(!\M_br_cond_taken_history[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_bht_ptr_nxt[1]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_bht_ptr_nxt[1] .extended_lut = "off";
defparam \F_bht_ptr_nxt[1] .lut_mask = 64'h6666666666666666;
defparam \F_bht_ptr_nxt[1] .shared_arith = "off";

dffeas \M_br_cond_taken_history[2] (
	.clk(clk_clk),
	.d(\M_br_cond_taken_history[1]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\M_br_cond_taken_history[0]~0_combout ),
	.q(\M_br_cond_taken_history[2]~q ),
	.prn(vcc));
defparam \M_br_cond_taken_history[2] .is_wysiwyg = "true";
defparam \M_br_cond_taken_history[2] .power_up = "low";

cyclonev_lcell_comb \F_bht_ptr_nxt[2] (
	.dataa(!\F_ic_data_rd_addr_nxt[2]~5_combout ),
	.datab(!\M_br_cond_taken_history[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_bht_ptr_nxt[2]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_bht_ptr_nxt[2] .extended_lut = "off";
defparam \F_bht_ptr_nxt[2] .lut_mask = 64'h6666666666666666;
defparam \F_bht_ptr_nxt[2] .shared_arith = "off";

dffeas \M_br_cond_taken_history[3] (
	.clk(clk_clk),
	.d(\M_br_cond_taken_history[2]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\M_br_cond_taken_history[0]~0_combout ),
	.q(\M_br_cond_taken_history[3]~q ),
	.prn(vcc));
defparam \M_br_cond_taken_history[3] .is_wysiwyg = "true";
defparam \M_br_cond_taken_history[3] .power_up = "low";

cyclonev_lcell_comb \F_bht_ptr_nxt[3] (
	.dataa(!\F_ic_tag_rd_addr_nxt[0]~5_combout ),
	.datab(!\M_br_cond_taken_history[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_bht_ptr_nxt[3]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_bht_ptr_nxt[3] .extended_lut = "off";
defparam \F_bht_ptr_nxt[3] .lut_mask = 64'h6666666666666666;
defparam \F_bht_ptr_nxt[3] .shared_arith = "off";

dffeas \M_br_cond_taken_history[4] (
	.clk(clk_clk),
	.d(\M_br_cond_taken_history[3]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\M_br_cond_taken_history[0]~0_combout ),
	.q(\M_br_cond_taken_history[4]~q ),
	.prn(vcc));
defparam \M_br_cond_taken_history[4] .is_wysiwyg = "true";
defparam \M_br_cond_taken_history[4] .power_up = "low";

cyclonev_lcell_comb \F_bht_ptr_nxt[4] (
	.dataa(!\F_ic_tag_rd_addr_nxt[1]~7_combout ),
	.datab(!\M_br_cond_taken_history[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_bht_ptr_nxt[4]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_bht_ptr_nxt[4] .extended_lut = "off";
defparam \F_bht_ptr_nxt[4] .lut_mask = 64'h6666666666666666;
defparam \F_bht_ptr_nxt[4] .shared_arith = "off";

dffeas \M_br_cond_taken_history[5] (
	.clk(clk_clk),
	.d(\M_br_cond_taken_history[4]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\M_br_cond_taken_history[0]~0_combout ),
	.q(\M_br_cond_taken_history[5]~q ),
	.prn(vcc));
defparam \M_br_cond_taken_history[5] .is_wysiwyg = "true";
defparam \M_br_cond_taken_history[5] .power_up = "low";

cyclonev_lcell_comb \F_bht_ptr_nxt[5] (
	.dataa(!\F_ic_tag_rd_addr_nxt[2]~9_combout ),
	.datab(!\M_br_cond_taken_history[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_bht_ptr_nxt[5]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_bht_ptr_nxt[5] .extended_lut = "off";
defparam \F_bht_ptr_nxt[5] .lut_mask = 64'h6666666666666666;
defparam \F_bht_ptr_nxt[5] .shared_arith = "off";

dffeas \M_br_cond_taken_history[6] (
	.clk(clk_clk),
	.d(\M_br_cond_taken_history[5]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\M_br_cond_taken_history[0]~0_combout ),
	.q(\M_br_cond_taken_history[6]~q ),
	.prn(vcc));
defparam \M_br_cond_taken_history[6] .is_wysiwyg = "true";
defparam \M_br_cond_taken_history[6] .power_up = "low";

cyclonev_lcell_comb \F_bht_ptr_nxt[6] (
	.dataa(!\F_ic_tag_rd_addr_nxt[3]~11_combout ),
	.datab(!\M_br_cond_taken_history[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_bht_ptr_nxt[6]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_bht_ptr_nxt[6] .extended_lut = "off";
defparam \F_bht_ptr_nxt[6] .lut_mask = 64'h6666666666666666;
defparam \F_bht_ptr_nxt[6] .shared_arith = "off";

dffeas \M_br_cond_taken_history[7] (
	.clk(clk_clk),
	.d(\M_br_cond_taken_history[6]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\M_br_cond_taken_history[0]~0_combout ),
	.q(\M_br_cond_taken_history[7]~q ),
	.prn(vcc));
defparam \M_br_cond_taken_history[7] .is_wysiwyg = "true";
defparam \M_br_cond_taken_history[7] .power_up = "low";

cyclonev_lcell_comb \F_bht_ptr_nxt[7] (
	.dataa(!\F_ic_tag_rd_addr_nxt[4]~13_combout ),
	.datab(!\M_br_cond_taken_history[7]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_bht_ptr_nxt[7]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_bht_ptr_nxt[7] .extended_lut = "off";
defparam \F_bht_ptr_nxt[7] .lut_mask = 64'h6666666666666666;
defparam \F_bht_ptr_nxt[7] .shared_arith = "off";

cyclonev_lcell_comb ic_tag_clr_valid_bits_nxt(
	.dataa(!clr_break_line1),
	.datab(!\A_valid_from_M~q ),
	.datac(!\D_ic_fill_starting~combout ),
	.datad(!\A_ctrl_invalidate_i~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_tag_clr_valid_bits_nxt~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam ic_tag_clr_valid_bits_nxt.extended_lut = "off";
defparam ic_tag_clr_valid_bits_nxt.lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam ic_tag_clr_valid_bits_nxt.shared_arith = "off";

cyclonev_lcell_comb \ic_tag_wraddress_nxt~6 (
	.dataa(!\A_valid_from_M~q ),
	.datab(!\A_inst_result[5]~q ),
	.datac(!\ic_tag_wraddress_nxt~0_combout ),
	.datad(!\A_ctrl_invalidate_i~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_tag_wraddress_nxt~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_tag_wraddress_nxt~6 .extended_lut = "off";
defparam \ic_tag_wraddress_nxt~6 .lut_mask = 64'h7FBF7FBF7FBF7FBF;
defparam \ic_tag_wraddress_nxt~6 .shared_arith = "off";

cyclonev_lcell_comb \ic_tag_wraddress_nxt[1]~7 (
	.dataa(!\A_valid_from_M~q ),
	.datab(!\A_inst_result[6]~q ),
	.datac(!\ic_tag_wraddress_nxt~5_combout ),
	.datad(!\A_ctrl_invalidate_i~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_tag_wraddress_nxt[1]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_tag_wraddress_nxt[1]~7 .extended_lut = "off";
defparam \ic_tag_wraddress_nxt[1]~7 .lut_mask = 64'h7FBF7FBF7FBF7FBF;
defparam \ic_tag_wraddress_nxt[1]~7 .shared_arith = "off";

cyclonev_lcell_comb \ic_tag_wraddress_nxt[2]~8 (
	.dataa(!\A_valid_from_M~q ),
	.datab(!\A_inst_result[7]~q ),
	.datac(!\ic_tag_wraddress_nxt~4_combout ),
	.datad(!\A_ctrl_invalidate_i~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_tag_wraddress_nxt[2]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_tag_wraddress_nxt[2]~8 .extended_lut = "off";
defparam \ic_tag_wraddress_nxt[2]~8 .lut_mask = 64'h7FBF7FBF7FBF7FBF;
defparam \ic_tag_wraddress_nxt[2]~8 .shared_arith = "off";

cyclonev_lcell_comb \ic_tag_wraddress_nxt[3]~9 (
	.dataa(!\A_valid_from_M~q ),
	.datab(!\A_inst_result[8]~q ),
	.datac(!\ic_tag_wraddress_nxt~3_combout ),
	.datad(!\A_ctrl_invalidate_i~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_tag_wraddress_nxt[3]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_tag_wraddress_nxt[3]~9 .extended_lut = "off";
defparam \ic_tag_wraddress_nxt[3]~9 .lut_mask = 64'h7FBF7FBF7FBF7FBF;
defparam \ic_tag_wraddress_nxt[3]~9 .shared_arith = "off";

cyclonev_lcell_comb \ic_tag_wraddress_nxt[4]~10 (
	.dataa(!\A_valid_from_M~q ),
	.datab(!\A_inst_result[9]~q ),
	.datac(!\ic_tag_wraddress_nxt~2_combout ),
	.datad(!\A_ctrl_invalidate_i~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_tag_wraddress_nxt[4]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_tag_wraddress_nxt[4]~10 .extended_lut = "off";
defparam \ic_tag_wraddress_nxt[4]~10 .lut_mask = 64'h7FBF7FBF7FBF7FBF;
defparam \ic_tag_wraddress_nxt[4]~10 .shared_arith = "off";

cyclonev_lcell_comb \ic_tag_wraddress_nxt[5]~11 (
	.dataa(!\A_valid_from_M~q ),
	.datab(!\A_inst_result[10]~q ),
	.datac(!\ic_tag_wraddress_nxt~1_combout ),
	.datad(!\A_ctrl_invalidate_i~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_tag_wraddress_nxt[5]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_tag_wraddress_nxt[5]~11 .extended_lut = "off";
defparam \ic_tag_wraddress_nxt[5]~11 .lut_mask = 64'h7FBF7FBF7FBF7FBF;
defparam \ic_tag_wraddress_nxt[5]~11 .shared_arith = "off";

dffeas \E_bht_data[0] (
	.clk(clk_clk),
	.d(\D_bht_data[0]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_bht_data[0]~q ),
	.prn(vcc));
defparam \E_bht_data[0] .is_wysiwyg = "true";
defparam \E_bht_data[0] .power_up = "low";

cyclonev_lcell_comb E_br_mispredict(
	.dataa(!\Add9~61_sumout ),
	.datab(!\E_br_result~0_combout ),
	.datac(!\E_br_result~1_combout ),
	.datad(!\E_bht_data[1]~q ),
	.datae(!\E_br_mispredict~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_br_mispredict~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam E_br_mispredict.extended_lut = "off";
defparam E_br_mispredict.lut_mask = 64'h6996FFFF6996FFFF;
defparam E_br_mispredict.shared_arith = "off";

dffeas \E_bht_ptr[0] (
	.clk(clk_clk),
	.d(\D_bht_ptr[0]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_bht_ptr[0]~q ),
	.prn(vcc));
defparam \E_bht_ptr[0] .is_wysiwyg = "true";
defparam \E_bht_ptr[0] .power_up = "low";

dffeas \E_bht_ptr[1] (
	.clk(clk_clk),
	.d(\D_bht_ptr[1]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_bht_ptr[1]~q ),
	.prn(vcc));
defparam \E_bht_ptr[1] .is_wysiwyg = "true";
defparam \E_bht_ptr[1] .power_up = "low";

dffeas \E_bht_ptr[2] (
	.clk(clk_clk),
	.d(\D_bht_ptr[2]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_bht_ptr[2]~q ),
	.prn(vcc));
defparam \E_bht_ptr[2] .is_wysiwyg = "true";
defparam \E_bht_ptr[2] .power_up = "low";

dffeas \E_bht_ptr[3] (
	.clk(clk_clk),
	.d(\D_bht_ptr[3]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_bht_ptr[3]~q ),
	.prn(vcc));
defparam \E_bht_ptr[3] .is_wysiwyg = "true";
defparam \E_bht_ptr[3] .power_up = "low";

dffeas \E_bht_ptr[4] (
	.clk(clk_clk),
	.d(\D_bht_ptr[4]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_bht_ptr[4]~q ),
	.prn(vcc));
defparam \E_bht_ptr[4] .is_wysiwyg = "true";
defparam \E_bht_ptr[4] .power_up = "low";

dffeas \E_bht_ptr[5] (
	.clk(clk_clk),
	.d(\D_bht_ptr[5]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_bht_ptr[5]~q ),
	.prn(vcc));
defparam \E_bht_ptr[5] .is_wysiwyg = "true";
defparam \E_bht_ptr[5] .power_up = "low";

dffeas \E_bht_ptr[6] (
	.clk(clk_clk),
	.d(\D_bht_ptr[6]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_bht_ptr[6]~q ),
	.prn(vcc));
defparam \E_bht_ptr[6] .is_wysiwyg = "true";
defparam \E_bht_ptr[6] .power_up = "low";

dffeas \E_bht_ptr[7] (
	.clk(clk_clk),
	.d(\D_bht_ptr[7]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_bht_ptr[7]~q ),
	.prn(vcc));
defparam \E_bht_ptr[7] .is_wysiwyg = "true";
defparam \E_bht_ptr[7] .power_up = "low";

cyclonev_lcell_comb \E_br_result~2 (
	.dataa(!\Add9~61_sumout ),
	.datab(!\E_br_result~0_combout ),
	.datac(!\E_br_result~1_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_br_result~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_br_result~2 .extended_lut = "off";
defparam \E_br_result~2 .lut_mask = 64'h2727272727272727;
defparam \E_br_result~2 .shared_arith = "off";

cyclonev_lcell_comb \M_br_cond_taken_history[0]~0 (
	.dataa(!\A_mem_stall~q ),
	.datab(!\E_br_mispredict~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_br_cond_taken_history[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_br_cond_taken_history[0]~0 .extended_lut = "off";
defparam \M_br_cond_taken_history[0]~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \M_br_cond_taken_history[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \ic_fill_valid_bits_nxt~0 (
	.dataa(!\D_ic_fill_starting_d1~q ),
	.datab(!\ic_fill_dp_offset_nxt[0]~1_combout ),
	.datac(!\ic_fill_dp_offset_nxt[1]~2_combout ),
	.datad(!\ic_fill_dp_offset_nxt[2]~0_combout ),
	.datae(!\ic_fill_valid_bits[5]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_valid_bits_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_valid_bits_nxt~0 .extended_lut = "off";
defparam \ic_fill_valid_bits_nxt~0 .lut_mask = 64'hFBFFFFFFFBFFFFFF;
defparam \ic_fill_valid_bits_nxt~0 .shared_arith = "off";

cyclonev_lcell_comb ic_fill_valid_bits_en(
	.dataa(!\ic_fill_dp_offset_en~0_combout ),
	.datab(!\ic_tag_clr_valid_bits_nxt~combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_valid_bits_en~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam ic_fill_valid_bits_en.extended_lut = "off";
defparam ic_fill_valid_bits_en.lut_mask = 64'h7777777777777777;
defparam ic_fill_valid_bits_en.shared_arith = "off";

cyclonev_lcell_comb \ic_fill_valid_bits_nxt~1 (
	.dataa(!\D_ic_fill_starting_d1~q ),
	.datab(!\ic_fill_dp_offset_nxt[0]~1_combout ),
	.datac(!\ic_fill_dp_offset_nxt[1]~2_combout ),
	.datad(!\ic_fill_dp_offset_nxt[2]~0_combout ),
	.datae(!\ic_fill_valid_bits[7]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_valid_bits_nxt~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_valid_bits_nxt~1 .extended_lut = "off";
defparam \ic_fill_valid_bits_nxt~1 .lut_mask = 64'hBFFFFFFFBFFFFFFF;
defparam \ic_fill_valid_bits_nxt~1 .shared_arith = "off";

cyclonev_lcell_comb \ic_fill_valid_bits_nxt~2 (
	.dataa(!\D_ic_fill_starting_d1~q ),
	.datab(!\ic_fill_dp_offset_nxt[0]~1_combout ),
	.datac(!\ic_fill_dp_offset_nxt[1]~2_combout ),
	.datad(!\ic_fill_dp_offset_nxt[2]~0_combout ),
	.datae(!\ic_fill_valid_bits[4]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_valid_bits_nxt~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_valid_bits_nxt~2 .extended_lut = "off";
defparam \ic_fill_valid_bits_nxt~2 .lut_mask = 64'hFEFFFFFFFEFFFFFF;
defparam \ic_fill_valid_bits_nxt~2 .shared_arith = "off";

cyclonev_lcell_comb \ic_fill_valid_bits_nxt~3 (
	.dataa(!\D_ic_fill_starting_d1~q ),
	.datab(!\ic_fill_dp_offset_nxt[0]~1_combout ),
	.datac(!\ic_fill_dp_offset_nxt[1]~2_combout ),
	.datad(!\ic_fill_dp_offset_nxt[2]~0_combout ),
	.datae(!\ic_fill_valid_bits[6]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_valid_bits_nxt~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_valid_bits_nxt~3 .extended_lut = "off";
defparam \ic_fill_valid_bits_nxt~3 .lut_mask = 64'hEFFFFFFFEFFFFFFF;
defparam \ic_fill_valid_bits_nxt~3 .shared_arith = "off";

dffeas \D_bht_data[0] (
	.clk(clk_clk),
	.d(\first_nios2_system_cpu_cpu_bht|the_altsyncram|auto_generated|q_b[0] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_bht_data[0]~q ),
	.prn(vcc));
defparam \D_bht_data[0] .is_wysiwyg = "true";
defparam \D_bht_data[0] .power_up = "low";

dffeas \D_bht_ptr[0] (
	.clk(clk_clk),
	.d(\F_bht_ptr[0]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_bht_ptr[0]~q ),
	.prn(vcc));
defparam \D_bht_ptr[0] .is_wysiwyg = "true";
defparam \D_bht_ptr[0] .power_up = "low";

dffeas \D_bht_ptr[1] (
	.clk(clk_clk),
	.d(\F_bht_ptr[1]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_bht_ptr[1]~q ),
	.prn(vcc));
defparam \D_bht_ptr[1] .is_wysiwyg = "true";
defparam \D_bht_ptr[1] .power_up = "low";

dffeas \D_bht_ptr[2] (
	.clk(clk_clk),
	.d(\F_bht_ptr[2]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_bht_ptr[2]~q ),
	.prn(vcc));
defparam \D_bht_ptr[2] .is_wysiwyg = "true";
defparam \D_bht_ptr[2] .power_up = "low";

dffeas \D_bht_ptr[3] (
	.clk(clk_clk),
	.d(\F_bht_ptr[3]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_bht_ptr[3]~q ),
	.prn(vcc));
defparam \D_bht_ptr[3] .is_wysiwyg = "true";
defparam \D_bht_ptr[3] .power_up = "low";

dffeas \D_bht_ptr[4] (
	.clk(clk_clk),
	.d(\F_bht_ptr[4]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_bht_ptr[4]~q ),
	.prn(vcc));
defparam \D_bht_ptr[4] .is_wysiwyg = "true";
defparam \D_bht_ptr[4] .power_up = "low";

dffeas \D_bht_ptr[5] (
	.clk(clk_clk),
	.d(\F_bht_ptr[5]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_bht_ptr[5]~q ),
	.prn(vcc));
defparam \D_bht_ptr[5] .is_wysiwyg = "true";
defparam \D_bht_ptr[5] .power_up = "low";

dffeas \D_bht_ptr[6] (
	.clk(clk_clk),
	.d(\F_bht_ptr[6]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_bht_ptr[6]~q ),
	.prn(vcc));
defparam \D_bht_ptr[6] .is_wysiwyg = "true";
defparam \D_bht_ptr[6] .power_up = "low";

dffeas \D_bht_ptr[7] (
	.clk(clk_clk),
	.d(\F_bht_ptr[7]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_bht_ptr[7]~q ),
	.prn(vcc));
defparam \D_bht_ptr[7] .is_wysiwyg = "true";
defparam \D_bht_ptr[7] .power_up = "low";

cyclonev_lcell_comb \ic_fill_valid_bits_nxt~4 (
	.dataa(!\D_ic_fill_starting_d1~q ),
	.datab(!\ic_fill_dp_offset_nxt[0]~1_combout ),
	.datac(!\ic_fill_dp_offset_nxt[1]~2_combout ),
	.datad(!\ic_fill_dp_offset_nxt[2]~0_combout ),
	.datae(!\ic_fill_valid_bits[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_valid_bits_nxt~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_valid_bits_nxt~4 .extended_lut = "off";
defparam \ic_fill_valid_bits_nxt~4 .lut_mask = 64'hFFFBFFFFFFFBFFFF;
defparam \ic_fill_valid_bits_nxt~4 .shared_arith = "off";

cyclonev_lcell_comb \ic_fill_valid_bits_nxt~5 (
	.dataa(!\D_ic_fill_starting_d1~q ),
	.datab(!\ic_fill_dp_offset_nxt[0]~1_combout ),
	.datac(!\ic_fill_dp_offset_nxt[1]~2_combout ),
	.datad(!\ic_fill_dp_offset_nxt[2]~0_combout ),
	.datae(!\ic_fill_valid_bits[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_valid_bits_nxt~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_valid_bits_nxt~5 .extended_lut = "off";
defparam \ic_fill_valid_bits_nxt~5 .lut_mask = 64'hFFBFFFFFFFBFFFFF;
defparam \ic_fill_valid_bits_nxt~5 .shared_arith = "off";

cyclonev_lcell_comb \ic_fill_valid_bits_nxt~6 (
	.dataa(!\D_ic_fill_starting_d1~q ),
	.datab(!\ic_fill_dp_offset_nxt[0]~1_combout ),
	.datac(!\ic_fill_dp_offset_nxt[1]~2_combout ),
	.datad(!\ic_fill_dp_offset_nxt[2]~0_combout ),
	.datae(!\ic_fill_valid_bits[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_valid_bits_nxt~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_valid_bits_nxt~6 .extended_lut = "off";
defparam \ic_fill_valid_bits_nxt~6 .lut_mask = 64'hFFFEFFFFFFFEFFFF;
defparam \ic_fill_valid_bits_nxt~6 .shared_arith = "off";

cyclonev_lcell_comb \ic_fill_valid_bits_nxt~7 (
	.dataa(!\D_ic_fill_starting_d1~q ),
	.datab(!\ic_fill_dp_offset_nxt[0]~1_combout ),
	.datac(!\ic_fill_dp_offset_nxt[1]~2_combout ),
	.datad(!\ic_fill_dp_offset_nxt[2]~0_combout ),
	.datae(!\ic_fill_valid_bits[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_valid_bits_nxt~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_valid_bits_nxt~7 .extended_lut = "off";
defparam \ic_fill_valid_bits_nxt~7 .lut_mask = 64'hFFEFFFFFFFEFFFFF;
defparam \ic_fill_valid_bits_nxt~7 .shared_arith = "off";

dffeas \F_bht_ptr[0] (
	.clk(clk_clk),
	.d(\F_bht_ptr_nxt[0]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\F_bht_ptr[0]~q ),
	.prn(vcc));
defparam \F_bht_ptr[0] .is_wysiwyg = "true";
defparam \F_bht_ptr[0] .power_up = "low";

dffeas \F_bht_ptr[1] (
	.clk(clk_clk),
	.d(\F_bht_ptr_nxt[1]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\F_bht_ptr[1]~q ),
	.prn(vcc));
defparam \F_bht_ptr[1] .is_wysiwyg = "true";
defparam \F_bht_ptr[1] .power_up = "low";

dffeas \F_bht_ptr[2] (
	.clk(clk_clk),
	.d(\F_bht_ptr_nxt[2]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\F_bht_ptr[2]~q ),
	.prn(vcc));
defparam \F_bht_ptr[2] .is_wysiwyg = "true";
defparam \F_bht_ptr[2] .power_up = "low";

dffeas \F_bht_ptr[3] (
	.clk(clk_clk),
	.d(\F_bht_ptr_nxt[3]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\F_bht_ptr[3]~q ),
	.prn(vcc));
defparam \F_bht_ptr[3] .is_wysiwyg = "true";
defparam \F_bht_ptr[3] .power_up = "low";

dffeas \F_bht_ptr[4] (
	.clk(clk_clk),
	.d(\F_bht_ptr_nxt[4]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\F_bht_ptr[4]~q ),
	.prn(vcc));
defparam \F_bht_ptr[4] .is_wysiwyg = "true";
defparam \F_bht_ptr[4] .power_up = "low";

dffeas \F_bht_ptr[5] (
	.clk(clk_clk),
	.d(\F_bht_ptr_nxt[5]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\F_bht_ptr[5]~q ),
	.prn(vcc));
defparam \F_bht_ptr[5] .is_wysiwyg = "true";
defparam \F_bht_ptr[5] .power_up = "low";

dffeas \F_bht_ptr[6] (
	.clk(clk_clk),
	.d(\F_bht_ptr_nxt[6]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\F_bht_ptr[6]~q ),
	.prn(vcc));
defparam \F_bht_ptr[6] .is_wysiwyg = "true";
defparam \F_bht_ptr[6] .power_up = "low";

dffeas \F_bht_ptr[7] (
	.clk(clk_clk),
	.d(\F_bht_ptr_nxt[7]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\F_bht_ptr[7]~q ),
	.prn(vcc));
defparam \F_bht_ptr[7] .is_wysiwyg = "true";
defparam \F_bht_ptr[7] .power_up = "low";

cyclonev_lcell_comb \ic_tag_clr_valid_bits~0 (
	.dataa(!\ic_tag_clr_valid_bits_nxt~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_tag_clr_valid_bits~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_tag_clr_valid_bits~0 .extended_lut = "off";
defparam \ic_tag_clr_valid_bits~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \ic_tag_clr_valid_bits~0 .shared_arith = "off";

cyclonev_lcell_comb \M_br_mispredict~_wirecell (
	.dataa(!\M_br_mispredict~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_br_mispredict~_wirecell_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_br_mispredict~_wirecell .extended_lut = "off";
defparam \M_br_mispredict~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \M_br_mispredict~_wirecell .shared_arith = "off";

dffeas \A_st_data[0] (
	.clk(clk_clk),
	.d(\M_st_data[0]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(A_st_data_0),
	.prn(vcc));
defparam \A_st_data[0] .is_wysiwyg = "true";
defparam \A_st_data[0] .power_up = "low";

dffeas \A_mem_baddr[4] (
	.clk(clk_clk),
	.d(\M_mem_baddr[4]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(A_mem_baddr_4),
	.prn(vcc));
defparam \A_mem_baddr[4] .is_wysiwyg = "true";
defparam \A_mem_baddr[4] .power_up = "low";

dffeas \A_mem_baddr[5] (
	.clk(clk_clk),
	.d(\M_mem_baddr[5]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(A_mem_baddr_5),
	.prn(vcc));
defparam \A_mem_baddr[5] .is_wysiwyg = "true";
defparam \A_mem_baddr[5] .power_up = "low";

dffeas \A_mem_baddr[8] (
	.clk(clk_clk),
	.d(\M_mem_baddr[8]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(A_mem_baddr_8),
	.prn(vcc));
defparam \A_mem_baddr[8] .is_wysiwyg = "true";
defparam \A_mem_baddr[8] .power_up = "low";

dffeas \A_mem_baddr[16] (
	.clk(clk_clk),
	.d(\M_mem_baddr[16]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(A_mem_baddr_16),
	.prn(vcc));
defparam \A_mem_baddr[16] .is_wysiwyg = "true";
defparam \A_mem_baddr[16] .power_up = "low";

dffeas \A_mem_baddr[15] (
	.clk(clk_clk),
	.d(\M_mem_baddr[15]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(A_mem_baddr_15),
	.prn(vcc));
defparam \A_mem_baddr[15] .is_wysiwyg = "true";
defparam \A_mem_baddr[15] .power_up = "low";

dffeas \A_mem_baddr[14] (
	.clk(clk_clk),
	.d(\M_mem_baddr[14]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(A_mem_baddr_14),
	.prn(vcc));
defparam \A_mem_baddr[14] .is_wysiwyg = "true";
defparam \A_mem_baddr[14] .power_up = "low";

dffeas \A_mem_baddr[13] (
	.clk(clk_clk),
	.d(\M_mem_baddr[13]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(A_mem_baddr_13),
	.prn(vcc));
defparam \A_mem_baddr[13] .is_wysiwyg = "true";
defparam \A_mem_baddr[13] .power_up = "low";

dffeas \A_mem_baddr[12] (
	.clk(clk_clk),
	.d(\M_mem_baddr[12]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(A_mem_baddr_12),
	.prn(vcc));
defparam \A_mem_baddr[12] .is_wysiwyg = "true";
defparam \A_mem_baddr[12] .power_up = "low";

dffeas \A_mem_baddr[11] (
	.clk(clk_clk),
	.d(\M_mem_baddr[11]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(A_mem_baddr_11),
	.prn(vcc));
defparam \A_mem_baddr[11] .is_wysiwyg = "true";
defparam \A_mem_baddr[11] .power_up = "low";

dffeas \A_mem_baddr[10] (
	.clk(clk_clk),
	.d(\M_mem_baddr[10]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(A_mem_baddr_10),
	.prn(vcc));
defparam \A_mem_baddr[10] .is_wysiwyg = "true";
defparam \A_mem_baddr[10] .power_up = "low";

dffeas \A_mem_baddr[9] (
	.clk(clk_clk),
	.d(\M_mem_baddr[9]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(A_mem_baddr_9),
	.prn(vcc));
defparam \A_mem_baddr[9] .is_wysiwyg = "true";
defparam \A_mem_baddr[9] .power_up = "low";

dffeas \A_mem_baddr[7] (
	.clk(clk_clk),
	.d(\M_mem_baddr[7]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(A_mem_baddr_7),
	.prn(vcc));
defparam \A_mem_baddr[7] .is_wysiwyg = "true";
defparam \A_mem_baddr[7] .power_up = "low";

dffeas \A_mem_baddr[6] (
	.clk(clk_clk),
	.d(\M_mem_baddr[6]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(A_mem_baddr_6),
	.prn(vcc));
defparam \A_mem_baddr[6] .is_wysiwyg = "true";
defparam \A_mem_baddr[6] .power_up = "low";

dffeas clr_break_line(
	.clk(clk_clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(clr_break_line1),
	.prn(vcc));
defparam clr_break_line.is_wysiwyg = "true";
defparam clr_break_line.power_up = "low";

dffeas d_write(
	.clk(clk_clk),
	.d(\d_write_nxt~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_write1),
	.prn(vcc));
defparam d_write.is_wysiwyg = "true";
defparam d_write.power_up = "low";

dffeas \A_mem_baddr[3] (
	.clk(clk_clk),
	.d(\M_mem_baddr[3]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(A_mem_baddr_3),
	.prn(vcc));
defparam \A_mem_baddr[3] .is_wysiwyg = "true";
defparam \A_mem_baddr[3] .power_up = "low";

dffeas \A_mem_baddr[2] (
	.clk(clk_clk),
	.d(\M_mem_baddr[2]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(A_mem_baddr_2),
	.prn(vcc));
defparam \A_mem_baddr[2] .is_wysiwyg = "true";
defparam \A_mem_baddr[2] .power_up = "low";

dffeas \A_st_data[1] (
	.clk(clk_clk),
	.d(\M_st_data[1]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(A_st_data_1),
	.prn(vcc));
defparam \A_st_data[1] .is_wysiwyg = "true";
defparam \A_st_data[1] .power_up = "low";

dffeas \A_st_data[2] (
	.clk(clk_clk),
	.d(\M_st_data[2]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(A_st_data_2),
	.prn(vcc));
defparam \A_st_data[2] .is_wysiwyg = "true";
defparam \A_st_data[2] .power_up = "low";

dffeas \A_st_data[3] (
	.clk(clk_clk),
	.d(\M_st_data[3]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(A_st_data_3),
	.prn(vcc));
defparam \A_st_data[3] .is_wysiwyg = "true";
defparam \A_st_data[3] .power_up = "low";

dffeas \A_st_data[4] (
	.clk(clk_clk),
	.d(\M_st_data[4]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(A_st_data_4),
	.prn(vcc));
defparam \A_st_data[4] .is_wysiwyg = "true";
defparam \A_st_data[4] .power_up = "low";

dffeas \A_st_data[5] (
	.clk(clk_clk),
	.d(\M_st_data[5]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(A_st_data_5),
	.prn(vcc));
defparam \A_st_data[5] .is_wysiwyg = "true";
defparam \A_st_data[5] .power_up = "low";

dffeas \A_st_data[6] (
	.clk(clk_clk),
	.d(\M_st_data[6]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(A_st_data_6),
	.prn(vcc));
defparam \A_st_data[6] .is_wysiwyg = "true";
defparam \A_st_data[6] .power_up = "low";

dffeas \A_st_data[7] (
	.clk(clk_clk),
	.d(\M_st_data[7]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(A_st_data_7),
	.prn(vcc));
defparam \A_st_data[7] .is_wysiwyg = "true";
defparam \A_st_data[7] .power_up = "low";

dffeas d_read(
	.clk(clk_clk),
	.d(\d_read_nxt~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_read1),
	.prn(vcc));
defparam d_read.is_wysiwyg = "true";
defparam d_read.power_up = "low";

dffeas W_debug_mode(
	.clk(clk_clk),
	.d(\W_debug_mode_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(W_debug_mode1),
	.prn(vcc));
defparam W_debug_mode.is_wysiwyg = "true";
defparam W_debug_mode.power_up = "low";

dffeas i_read(
	.clk(clk_clk),
	.d(\i_read_nxt~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(i_read1),
	.prn(vcc));
defparam i_read.is_wysiwyg = "true";
defparam i_read.power_up = "low";

dffeas \ic_fill_tag[5] (
	.clk(clk_clk),
	.d(\D_pc[14]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\D_ic_fill_starting~combout ),
	.q(ic_fill_tag_5),
	.prn(vcc));
defparam \ic_fill_tag[5] .is_wysiwyg = "true";
defparam \ic_fill_tag[5] .power_up = "low";

dffeas \ic_fill_tag[4] (
	.clk(clk_clk),
	.d(\D_pc[13]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\D_ic_fill_starting~combout ),
	.q(ic_fill_tag_4),
	.prn(vcc));
defparam \ic_fill_tag[4] .is_wysiwyg = "true";
defparam \ic_fill_tag[4] .power_up = "low";

dffeas \ic_fill_tag[3] (
	.clk(clk_clk),
	.d(\D_pc[12]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\D_ic_fill_starting~combout ),
	.q(ic_fill_tag_3),
	.prn(vcc));
defparam \ic_fill_tag[3] .is_wysiwyg = "true";
defparam \ic_fill_tag[3] .power_up = "low";

dffeas \ic_fill_tag[2] (
	.clk(clk_clk),
	.d(\D_pc[11]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\D_ic_fill_starting~combout ),
	.q(ic_fill_tag_2),
	.prn(vcc));
defparam \ic_fill_tag[2] .is_wysiwyg = "true";
defparam \ic_fill_tag[2] .power_up = "low";

dffeas \ic_fill_tag[1] (
	.clk(clk_clk),
	.d(\D_pc[10]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\D_ic_fill_starting~combout ),
	.q(ic_fill_tag_1),
	.prn(vcc));
defparam \ic_fill_tag[1] .is_wysiwyg = "true";
defparam \ic_fill_tag[1] .power_up = "low";

dffeas \ic_fill_tag[0] (
	.clk(clk_clk),
	.d(\D_pc[9]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\D_ic_fill_starting~combout ),
	.q(ic_fill_tag_0),
	.prn(vcc));
defparam \ic_fill_tag[0] .is_wysiwyg = "true";
defparam \ic_fill_tag[0] .power_up = "low";

dffeas \ic_fill_ap_offset[0] (
	.clk(clk_clk),
	.d(\ic_fill_ap_offset_nxt[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ic_fill_ap_offset[2]~0_combout ),
	.q(ic_fill_ap_offset_0),
	.prn(vcc));
defparam \ic_fill_ap_offset[0] .is_wysiwyg = "true";
defparam \ic_fill_ap_offset[0] .power_up = "low";

dffeas \ic_fill_line[0] (
	.clk(clk_clk),
	.d(\ic_tag_wraddress_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ic_fill_line_0),
	.prn(vcc));
defparam \ic_fill_line[0] .is_wysiwyg = "true";
defparam \ic_fill_line[0] .power_up = "low";

dffeas \ic_fill_ap_offset[2] (
	.clk(clk_clk),
	.d(\ic_fill_ap_offset_nxt[2]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ic_fill_ap_offset[2]~0_combout ),
	.q(ic_fill_ap_offset_2),
	.prn(vcc));
defparam \ic_fill_ap_offset[2] .is_wysiwyg = "true";
defparam \ic_fill_ap_offset[2] .power_up = "low";

dffeas \ic_fill_ap_offset[1] (
	.clk(clk_clk),
	.d(\ic_fill_ap_offset_nxt[1]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ic_fill_ap_offset[2]~0_combout ),
	.q(ic_fill_ap_offset_1),
	.prn(vcc));
defparam \ic_fill_ap_offset[1] .is_wysiwyg = "true";
defparam \ic_fill_ap_offset[1] .power_up = "low";

dffeas \ic_fill_line[5] (
	.clk(clk_clk),
	.d(\ic_tag_wraddress_nxt~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ic_fill_line_5),
	.prn(vcc));
defparam \ic_fill_line[5] .is_wysiwyg = "true";
defparam \ic_fill_line[5] .power_up = "low";

dffeas \ic_fill_line[4] (
	.clk(clk_clk),
	.d(\ic_tag_wraddress_nxt~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ic_fill_line_4),
	.prn(vcc));
defparam \ic_fill_line[4] .is_wysiwyg = "true";
defparam \ic_fill_line[4] .power_up = "low";

dffeas \ic_fill_line[3] (
	.clk(clk_clk),
	.d(\ic_tag_wraddress_nxt~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ic_fill_line_3),
	.prn(vcc));
defparam \ic_fill_line[3] .is_wysiwyg = "true";
defparam \ic_fill_line[3] .power_up = "low";

dffeas \ic_fill_line[2] (
	.clk(clk_clk),
	.d(\ic_tag_wraddress_nxt~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ic_fill_line_2),
	.prn(vcc));
defparam \ic_fill_line[2] .is_wysiwyg = "true";
defparam \ic_fill_line[2] .power_up = "low";

dffeas \ic_fill_line[1] (
	.clk(clk_clk),
	.d(\ic_tag_wraddress_nxt~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ic_fill_line_1),
	.prn(vcc));
defparam \ic_fill_line[1] .is_wysiwyg = "true";
defparam \ic_fill_line[1] .power_up = "low";

dffeas \A_mem_byte_en[0] (
	.clk(clk_clk),
	.d(\M_mem_byte_en[0]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(A_mem_byte_en_0),
	.prn(vcc));
defparam \A_mem_byte_en[0] .is_wysiwyg = "true";
defparam \A_mem_byte_en[0] .power_up = "low";

dffeas \A_st_data[16] (
	.clk(clk_clk),
	.d(\M_st_data[16]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(A_st_data_16),
	.prn(vcc));
defparam \A_st_data[16] .is_wysiwyg = "true";
defparam \A_st_data[16] .power_up = "low";

dffeas \A_st_data[22] (
	.clk(clk_clk),
	.d(\M_st_data[22]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(A_st_data_22),
	.prn(vcc));
defparam \A_st_data[22] .is_wysiwyg = "true";
defparam \A_st_data[22] .power_up = "low";

dffeas \A_mem_byte_en[2] (
	.clk(clk_clk),
	.d(\M_mem_byte_en[2]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(A_mem_byte_en_2),
	.prn(vcc));
defparam \A_mem_byte_en[2] .is_wysiwyg = "true";
defparam \A_mem_byte_en[2] .power_up = "low";

dffeas \A_st_data[23] (
	.clk(clk_clk),
	.d(\M_st_data[23]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(A_st_data_23),
	.prn(vcc));
defparam \A_st_data[23] .is_wysiwyg = "true";
defparam \A_st_data[23] .power_up = "low";

dffeas \A_st_data[24] (
	.clk(clk_clk),
	.d(\M_st_data[24]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(A_st_data_24),
	.prn(vcc));
defparam \A_st_data[24] .is_wysiwyg = "true";
defparam \A_st_data[24] .power_up = "low";

dffeas \A_mem_byte_en[3] (
	.clk(clk_clk),
	.d(\M_mem_byte_en[3]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(A_mem_byte_en_3),
	.prn(vcc));
defparam \A_mem_byte_en[3] .is_wysiwyg = "true";
defparam \A_mem_byte_en[3] .power_up = "low";

dffeas \A_st_data[25] (
	.clk(clk_clk),
	.d(\M_st_data[25]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(A_st_data_25),
	.prn(vcc));
defparam \A_st_data[25] .is_wysiwyg = "true";
defparam \A_st_data[25] .power_up = "low";

dffeas \A_st_data[31] (
	.clk(clk_clk),
	.d(\M_st_data[31]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(A_st_data_31),
	.prn(vcc));
defparam \A_st_data[31] .is_wysiwyg = "true";
defparam \A_st_data[31] .power_up = "low";

dffeas \A_st_data[21] (
	.clk(clk_clk),
	.d(\M_st_data[21]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(A_st_data_21),
	.prn(vcc));
defparam \A_st_data[21] .is_wysiwyg = "true";
defparam \A_st_data[21] .power_up = "low";

dffeas \A_st_data[11] (
	.clk(clk_clk),
	.d(\M_st_data[11]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(A_st_data_11),
	.prn(vcc));
defparam \A_st_data[11] .is_wysiwyg = "true";
defparam \A_st_data[11] .power_up = "low";

dffeas \A_mem_byte_en[1] (
	.clk(clk_clk),
	.d(\M_mem_byte_en[1]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(A_mem_byte_en_1),
	.prn(vcc));
defparam \A_mem_byte_en[1] .is_wysiwyg = "true";
defparam \A_mem_byte_en[1] .power_up = "low";

dffeas \A_st_data[28] (
	.clk(clk_clk),
	.d(\M_st_data[28]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(A_st_data_28),
	.prn(vcc));
defparam \A_st_data[28] .is_wysiwyg = "true";
defparam \A_st_data[28] .power_up = "low";

dffeas \A_st_data[10] (
	.clk(clk_clk),
	.d(\M_st_data[10]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(A_st_data_10),
	.prn(vcc));
defparam \A_st_data[10] .is_wysiwyg = "true";
defparam \A_st_data[10] .power_up = "low";

dffeas \A_st_data[27] (
	.clk(clk_clk),
	.d(\M_st_data[27]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(A_st_data_27),
	.prn(vcc));
defparam \A_st_data[27] .is_wysiwyg = "true";
defparam \A_st_data[27] .power_up = "low";

dffeas \A_st_data[8] (
	.clk(clk_clk),
	.d(\M_st_data[8]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(A_st_data_8),
	.prn(vcc));
defparam \A_st_data[8] .is_wysiwyg = "true";
defparam \A_st_data[8] .power_up = "low";

dffeas \A_st_data[9] (
	.clk(clk_clk),
	.d(\M_st_data[9]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(A_st_data_9),
	.prn(vcc));
defparam \A_st_data[9] .is_wysiwyg = "true";
defparam \A_st_data[9] .power_up = "low";

dffeas \A_st_data[26] (
	.clk(clk_clk),
	.d(\M_st_data[26]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(A_st_data_26),
	.prn(vcc));
defparam \A_st_data[26] .is_wysiwyg = "true";
defparam \A_st_data[26] .power_up = "low";

dffeas \A_st_data[20] (
	.clk(clk_clk),
	.d(\M_st_data[20]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(A_st_data_20),
	.prn(vcc));
defparam \A_st_data[20] .is_wysiwyg = "true";
defparam \A_st_data[20] .power_up = "low";

dffeas \A_st_data[19] (
	.clk(clk_clk),
	.d(\M_st_data[19]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(A_st_data_19),
	.prn(vcc));
defparam \A_st_data[19] .is_wysiwyg = "true";
defparam \A_st_data[19] .power_up = "low";

dffeas \A_st_data[17] (
	.clk(clk_clk),
	.d(\M_st_data[17]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(A_st_data_17),
	.prn(vcc));
defparam \A_st_data[17] .is_wysiwyg = "true";
defparam \A_st_data[17] .power_up = "low";

dffeas \A_st_data[30] (
	.clk(clk_clk),
	.d(\M_st_data[30]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(A_st_data_30),
	.prn(vcc));
defparam \A_st_data[30] .is_wysiwyg = "true";
defparam \A_st_data[30] .power_up = "low";

dffeas \A_st_data[18] (
	.clk(clk_clk),
	.d(\M_st_data[18]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(A_st_data_18),
	.prn(vcc));
defparam \A_st_data[18] .is_wysiwyg = "true";
defparam \A_st_data[18] .power_up = "low";

dffeas \A_st_data[15] (
	.clk(clk_clk),
	.d(\M_st_data[15]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(A_st_data_15),
	.prn(vcc));
defparam \A_st_data[15] .is_wysiwyg = "true";
defparam \A_st_data[15] .power_up = "low";

dffeas \A_st_data[12] (
	.clk(clk_clk),
	.d(\M_st_data[12]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(A_st_data_12),
	.prn(vcc));
defparam \A_st_data[12] .is_wysiwyg = "true";
defparam \A_st_data[12] .power_up = "low";

dffeas \A_st_data[13] (
	.clk(clk_clk),
	.d(\M_st_data[13]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(A_st_data_13),
	.prn(vcc));
defparam \A_st_data[13] .is_wysiwyg = "true";
defparam \A_st_data[13] .power_up = "low";

dffeas \A_st_data[14] (
	.clk(clk_clk),
	.d(\M_st_data[14]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(A_st_data_14),
	.prn(vcc));
defparam \A_st_data[14] .is_wysiwyg = "true";
defparam \A_st_data[14] .power_up = "low";

dffeas \A_st_data[29] (
	.clk(clk_clk),
	.d(\M_st_data[29]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(A_st_data_29),
	.prn(vcc));
defparam \A_st_data[29] .is_wysiwyg = "true";
defparam \A_st_data[29] .power_up = "low";

dffeas M_sel_data_master(
	.clk(clk_clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_sel_data_master~q ),
	.prn(vcc));
defparam M_sel_data_master.is_wysiwyg = "true";
defparam M_sel_data_master.power_up = "low";

dffeas A_valid_from_M(
	.clk(clk_clk),
	.d(\M_valid~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_valid_from_M~q ),
	.prn(vcc));
defparam A_valid_from_M.is_wysiwyg = "true";
defparam A_valid_from_M.power_up = "low";

dffeas \D_iw[0] (
	.clk(clk_clk),
	.d(\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[0] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_iw[0]~q ),
	.prn(vcc));
defparam \D_iw[0] .is_wysiwyg = "true";
defparam \D_iw[0] .power_up = "low";

dffeas \D_iw[1] (
	.clk(clk_clk),
	.d(\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[1] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_iw[1]~q ),
	.prn(vcc));
defparam \D_iw[1] .is_wysiwyg = "true";
defparam \D_iw[1] .power_up = "low";

dffeas \D_iw[2] (
	.clk(clk_clk),
	.d(\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[2] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_iw[2]~q ),
	.prn(vcc));
defparam \D_iw[2] .is_wysiwyg = "true";
defparam \D_iw[2] .power_up = "low";

dffeas \D_iw[3] (
	.clk(clk_clk),
	.d(\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[3] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_iw[3]~q ),
	.prn(vcc));
defparam \D_iw[3] .is_wysiwyg = "true";
defparam \D_iw[3] .power_up = "low";

dffeas \D_iw[4] (
	.clk(clk_clk),
	.d(\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[4] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_iw[4]~q ),
	.prn(vcc));
defparam \D_iw[4] .is_wysiwyg = "true";
defparam \D_iw[4] .power_up = "low";

cyclonev_lcell_comb \Equal95~0 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[1]~q ),
	.datac(!\D_iw[2]~q ),
	.datad(!\D_iw[3]~q ),
	.datae(!\D_iw[4]~q ),
	.dataf(!\D_iw[5]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal95~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal95~0 .extended_lut = "off";
defparam \Equal95~0 .lut_mask = 64'hFBFFFFFFFFFFFFFF;
defparam \Equal95~0 .shared_arith = "off";

dffeas \D_iw[16] (
	.clk(clk_clk),
	.d(\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[16] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_iw[16]~q ),
	.prn(vcc));
defparam \D_iw[16] .is_wysiwyg = "true";
defparam \D_iw[16] .power_up = "low";

dffeas \D_iw[15] (
	.clk(clk_clk),
	.d(\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[15] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_iw[15]~q ),
	.prn(vcc));
defparam \D_iw[15] .is_wysiwyg = "true";
defparam \D_iw[15] .power_up = "low";

dffeas \D_iw[14] (
	.clk(clk_clk),
	.d(\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[14] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_iw[14]~q ),
	.prn(vcc));
defparam \D_iw[14] .is_wysiwyg = "true";
defparam \D_iw[14] .power_up = "low";

dffeas \D_iw[13] (
	.clk(clk_clk),
	.d(\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[13] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_iw[13]~q ),
	.prn(vcc));
defparam \D_iw[13] .is_wysiwyg = "true";
defparam \D_iw[13] .power_up = "low";

dffeas \D_iw[12] (
	.clk(clk_clk),
	.d(\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[12] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_iw[12]~q ),
	.prn(vcc));
defparam \D_iw[12] .is_wysiwyg = "true";
defparam \D_iw[12] .power_up = "low";

dffeas \D_iw[11] (
	.clk(clk_clk),
	.d(\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[11] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_iw[11]~q ),
	.prn(vcc));
defparam \D_iw[11] .is_wysiwyg = "true";
defparam \D_iw[11] .power_up = "low";

cyclonev_lcell_comb \D_ctrl_shift_rot~2 (
	.dataa(!\D_iw[16]~q ),
	.datab(!\D_iw[15]~q ),
	.datac(!\D_iw[14]~q ),
	.datad(!\D_iw[13]~q ),
	.datae(!\D_iw[12]~q ),
	.dataf(!\D_iw[11]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_shift_rot~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_shift_rot~2 .extended_lut = "off";
defparam \D_ctrl_shift_rot~2 .lut_mask = 64'hFFFFFFFFFFDFFFFF;
defparam \D_ctrl_shift_rot~2 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_late_result~3 (
	.dataa(!\D_iw[16]~q ),
	.datab(!\D_iw[14]~q ),
	.datac(!\D_iw[13]~q ),
	.datad(!\D_iw[12]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_late_result~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_late_result~3 .extended_lut = "off";
defparam \D_ctrl_late_result~3 .lut_mask = 64'hFDFFFDFFFDFFFDFF;
defparam \D_ctrl_late_result~3 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_illegal~4 (
	.dataa(!\D_iw[16]~q ),
	.datab(!\D_iw[15]~q ),
	.datac(!\D_iw[14]~q ),
	.datad(!\D_iw[13]~q ),
	.datae(!\D_iw[12]~q ),
	.dataf(!\D_iw[11]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_illegal~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_illegal~4 .extended_lut = "off";
defparam \D_ctrl_illegal~4 .lut_mask = 64'h6996966996696996;
defparam \D_ctrl_illegal~4 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_illegal~2 (
	.dataa(!\D_ctrl_shift_rot~2_combout ),
	.datab(!\D_ctrl_late_result~3_combout ),
	.datac(!\D_ctrl_illegal~4_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_illegal~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_illegal~2 .extended_lut = "off";
defparam \D_ctrl_illegal~2 .lut_mask = 64'hFEFEFEFEFEFEFEFE;
defparam \D_ctrl_illegal~2 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_flush_pipe_always~2 (
	.dataa(!\D_iw[5]~q ),
	.datab(!\D_iw[4]~q ),
	.datac(!\D_iw[3]~q ),
	.datad(!\D_iw[2]~q ),
	.datae(!\D_iw[1]~q ),
	.dataf(!\D_iw[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_flush_pipe_always~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_flush_pipe_always~2 .extended_lut = "off";
defparam \D_ctrl_flush_pipe_always~2 .lut_mask = 64'h9F6F6F9F6F9F9F6F;
defparam \D_ctrl_flush_pipe_always~2 .shared_arith = "off";

cyclonev_lcell_comb \Equal149~6 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[13]~q ),
	.datad(!\D_iw[14]~q ),
	.datae(!\D_iw[15]~q ),
	.dataf(!\D_iw[16]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal149~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal149~6 .extended_lut = "off";
defparam \Equal149~6 .lut_mask = 64'hFFEFFFFFFFFFFFFF;
defparam \Equal149~6 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_flush_pipe_always~0 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[13]~q ),
	.datad(!\D_iw[14]~q ),
	.datae(!\D_iw[15]~q ),
	.dataf(!\D_iw[16]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_flush_pipe_always~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_flush_pipe_always~0 .extended_lut = "off";
defparam \D_ctrl_flush_pipe_always~0 .lut_mask = 64'h6996966996696996;
defparam \D_ctrl_flush_pipe_always~0 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_flush_pipe_always~1 (
	.dataa(!\Equal95~0_combout ),
	.datab(!\D_ctrl_illegal~2_combout ),
	.datac(!\D_ctrl_flush_pipe_always~2_combout ),
	.datad(!\Equal149~6_combout ),
	.datae(!\D_ctrl_flush_pipe_always~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_flush_pipe_always~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_flush_pipe_always~1 .extended_lut = "off";
defparam \D_ctrl_flush_pipe_always~1 .lut_mask = 64'hDFFFFFFFDFFFFFFF;
defparam \D_ctrl_flush_pipe_always~1 .shared_arith = "off";

dffeas E_ctrl_flush_pipe_always(
	.clk(clk_clk),
	.d(\D_ctrl_flush_pipe_always~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_ctrl_flush_pipe_always~q ),
	.prn(vcc));
defparam E_ctrl_flush_pipe_always.is_wysiwyg = "true";
defparam E_ctrl_flush_pipe_always.power_up = "low";

dffeas M_ctrl_flush_pipe_always(
	.clk(clk_clk),
	.d(\E_ctrl_flush_pipe_always~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_ctrl_flush_pipe_always~q ),
	.prn(vcc));
defparam M_ctrl_flush_pipe_always.is_wysiwyg = "true";
defparam M_ctrl_flush_pipe_always.power_up = "low";

cyclonev_lcell_comb \A_pipe_flush_nxt~0 (
	.dataa(!\M_exc_allowed~0_combout ),
	.datab(!\M_exc_any~combout ),
	.datac(!\M_ctrl_flush_pipe_always~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_pipe_flush_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_pipe_flush_nxt~0 .extended_lut = "off";
defparam \A_pipe_flush_nxt~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \A_pipe_flush_nxt~0 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_cmp~4 (
	.dataa(!\D_iw[15]~q ),
	.datab(!\D_iw[14]~q ),
	.datac(!\D_iw[13]~q ),
	.datad(!\D_iw[12]~q ),
	.datae(!\D_iw[11]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_cmp~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_cmp~4 .extended_lut = "off";
defparam \D_ctrl_cmp~4 .lut_mask = 64'hFFFFFFF6FFFFFFF6;
defparam \D_ctrl_cmp~4 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_alu_force_xor~3 (
	.dataa(!\D_iw[4]~q ),
	.datab(!\D_iw[3]~q ),
	.datac(!\D_iw[2]~q ),
	.datad(!\D_iw[1]~q ),
	.datae(!\D_iw[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_alu_force_xor~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_alu_force_xor~3 .extended_lut = "off";
defparam \D_ctrl_alu_force_xor~3 .lut_mask = 64'hFFFFFBFFFFFFFBFF;
defparam \D_ctrl_alu_force_xor~3 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_alu_subtract~0 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[13]~q ),
	.datad(!\D_iw[14]~q ),
	.datae(!\D_iw[15]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_alu_subtract~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_alu_subtract~0 .extended_lut = "off";
defparam \D_ctrl_alu_subtract~0 .lut_mask = 64'hFDFFFFFFFDFFFFFF;
defparam \D_ctrl_alu_subtract~0 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_alu_subtract~2 (
	.dataa(!\D_iw[4]~q ),
	.datab(!\D_iw[3]~q ),
	.datac(!\D_iw[2]~q ),
	.datad(!\D_iw[1]~q ),
	.datae(!\D_iw[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_alu_subtract~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_alu_subtract~2 .extended_lut = "off";
defparam \D_ctrl_alu_subtract~2 .lut_mask = 64'hFFFFDFFDFFFFDFFD;
defparam \D_ctrl_alu_subtract~2 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_alu_subtract~1 (
	.dataa(!\Equal95~0_combout ),
	.datab(!\D_ctrl_cmp~4_combout ),
	.datac(!\D_ctrl_alu_force_xor~3_combout ),
	.datad(!\D_ctrl_alu_subtract~0_combout ),
	.datae(!\D_ctrl_alu_subtract~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_alu_subtract~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_alu_subtract~1 .extended_lut = "off";
defparam \D_ctrl_alu_subtract~1 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \D_ctrl_alu_subtract~1 .shared_arith = "off";

dffeas E_ctrl_alu_subtract(
	.clk(clk_clk),
	.d(\D_ctrl_alu_subtract~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_ctrl_alu_subtract~q ),
	.prn(vcc));
defparam E_ctrl_alu_subtract.is_wysiwyg = "true";
defparam E_ctrl_alu_subtract.power_up = "low";

cyclonev_lcell_comb \Equal149~3 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[13]~q ),
	.datad(!\D_iw[14]~q ),
	.datae(!\D_iw[15]~q ),
	.dataf(!\D_iw[16]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal149~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal149~3 .extended_lut = "off";
defparam \Equal149~3 .lut_mask = 64'hFFFFFFFFFFFEFFFF;
defparam \Equal149~3 .shared_arith = "off";

cyclonev_lcell_comb \Equal149~4 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[13]~q ),
	.datad(!\D_iw[14]~q ),
	.datae(!\D_iw[15]~q ),
	.dataf(!\D_iw[16]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal149~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal149~4 .extended_lut = "off";
defparam \Equal149~4 .lut_mask = 64'hFFFFFFFFFFFFFEFF;
defparam \Equal149~4 .shared_arith = "off";

cyclonev_lcell_comb \Equal95~1 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[1]~q ),
	.datac(!\D_iw[2]~q ),
	.datad(!\D_iw[3]~q ),
	.datae(!\D_iw[4]~q ),
	.dataf(!\D_iw[5]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal95~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal95~1 .extended_lut = "off";
defparam \Equal95~1 .lut_mask = 64'hFFFFFFFFFFFFFEFF;
defparam \Equal95~1 .shared_arith = "off";

cyclonev_lcell_comb \Equal95~2 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[1]~q ),
	.datac(!\D_iw[2]~q ),
	.datad(!\D_iw[3]~q ),
	.datae(!\D_iw[4]~q ),
	.dataf(!\D_iw[5]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal95~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal95~2 .extended_lut = "off";
defparam \Equal95~2 .lut_mask = 64'hFFFFFFFFFFFEFFFF;
defparam \Equal95~2 .shared_arith = "off";

cyclonev_lcell_comb \Equal95~3 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[1]~q ),
	.datac(!\D_iw[2]~q ),
	.datad(!\D_iw[3]~q ),
	.datae(!\D_iw[4]~q ),
	.dataf(!\D_iw[5]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal95~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal95~3 .extended_lut = "off";
defparam \Equal95~3 .lut_mask = 64'hFFFFFFFFFFFFBFFF;
defparam \Equal95~3 .shared_arith = "off";

cyclonev_lcell_comb \Equal95~5 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[1]~q ),
	.datac(!\D_iw[2]~q ),
	.datad(!\D_iw[3]~q ),
	.datae(!\D_iw[4]~q ),
	.dataf(!\D_iw[5]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal95~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal95~5 .extended_lut = "off";
defparam \Equal95~5 .lut_mask = 64'hFFFFFFFFFFBFFFFF;
defparam \Equal95~5 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_alu_signed_comparison~0 (
	.dataa(!\Equal95~1_combout ),
	.datab(!\Equal95~2_combout ),
	.datac(!\Equal95~3_combout ),
	.datad(!\Equal95~5_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_alu_signed_comparison~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_alu_signed_comparison~0 .extended_lut = "off";
defparam \D_ctrl_alu_signed_comparison~0 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \D_ctrl_alu_signed_comparison~0 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_alu_signed_comparison~1 (
	.dataa(!\Equal95~0_combout ),
	.datab(!\Equal149~3_combout ),
	.datac(!\Equal149~4_combout ),
	.datad(!\D_ctrl_alu_signed_comparison~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_alu_signed_comparison~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_alu_signed_comparison~1 .extended_lut = "off";
defparam \D_ctrl_alu_signed_comparison~1 .lut_mask = 64'hFF7FFF7FFF7FFF7F;
defparam \D_ctrl_alu_signed_comparison~1 .shared_arith = "off";

dffeas E_ctrl_alu_signed_comparison(
	.clk(clk_clk),
	.d(\D_ctrl_alu_signed_comparison~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_ctrl_alu_signed_comparison~q ),
	.prn(vcc));
defparam E_ctrl_alu_signed_comparison.is_wysiwyg = "true";
defparam E_ctrl_alu_signed_comparison.power_up = "low";

dffeas \D_iw[26] (
	.clk(clk_clk),
	.d(\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[26] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_iw[26]~q ),
	.prn(vcc));
defparam \D_iw[26] .is_wysiwyg = "true";
defparam \D_iw[26] .power_up = "low";

dffeas \D_iw[25] (
	.clk(clk_clk),
	.d(\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[25] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_iw[25]~q ),
	.prn(vcc));
defparam \D_iw[25] .is_wysiwyg = "true";
defparam \D_iw[25] .power_up = "low";

dffeas \D_iw[24] (
	.clk(clk_clk),
	.d(\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[24] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_iw[24]~q ),
	.prn(vcc));
defparam \D_iw[24] .is_wysiwyg = "true";
defparam \D_iw[24] .power_up = "low";

dffeas \D_iw[23] (
	.clk(clk_clk),
	.d(\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[23] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_iw[23]~q ),
	.prn(vcc));
defparam \D_iw[23] .is_wysiwyg = "true";
defparam \D_iw[23] .power_up = "low";

dffeas \D_iw[22] (
	.clk(clk_clk),
	.d(\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[22] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_iw[22]~q ),
	.prn(vcc));
defparam \D_iw[22] .is_wysiwyg = "true";
defparam \D_iw[22] .power_up = "low";

cyclonev_lcell_comb \Equal304~0 (
	.dataa(!\D_iw[26]~q ),
	.datab(!\D_iw[25]~q ),
	.datac(!\D_iw[24]~q ),
	.datad(!\D_iw[23]~q ),
	.datae(!\D_iw[22]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal304~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal304~0 .extended_lut = "off";
defparam \Equal304~0 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \Equal304~0 .shared_arith = "off";

cyclonev_lcell_comb \F_ctrl_b_is_dst~0 (
	.dataa(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[1] ),
	.datab(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[0] ),
	.datac(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[2] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ctrl_b_is_dst~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ctrl_b_is_dst~0 .extended_lut = "off";
defparam \F_ctrl_b_is_dst~0 .lut_mask = 64'hF6F6F6F6F6F6F6F6;
defparam \F_ctrl_b_is_dst~0 .shared_arith = "off";

dffeas D_ctrl_b_is_dst(
	.clk(clk_clk),
	.d(\F_ctrl_b_is_dst~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_ctrl_b_is_dst~q ),
	.prn(vcc));
defparam D_ctrl_b_is_dst.is_wysiwyg = "true";
defparam D_ctrl_b_is_dst.power_up = "low";

dffeas \D_iw[18] (
	.clk(clk_clk),
	.d(\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[18] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_iw[18]~q ),
	.prn(vcc));
defparam \D_iw[18] .is_wysiwyg = "true";
defparam \D_iw[18] .power_up = "low";

cyclonev_lcell_comb \F_ctrl_implicit_dst_retaddr~0 (
	.dataa(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[0] ),
	.datab(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[2] ),
	.datac(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[3] ),
	.datad(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[4] ),
	.datae(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[5] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ctrl_implicit_dst_retaddr~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ctrl_implicit_dst_retaddr~0 .extended_lut = "off";
defparam \F_ctrl_implicit_dst_retaddr~0 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \F_ctrl_implicit_dst_retaddr~0 .shared_arith = "off";

dffeas D_ctrl_implicit_dst_retaddr(
	.clk(clk_clk),
	.d(\F_ctrl_implicit_dst_retaddr~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_ctrl_implicit_dst_retaddr~q ),
	.prn(vcc));
defparam D_ctrl_implicit_dst_retaddr.is_wysiwyg = "true";
defparam D_ctrl_implicit_dst_retaddr.power_up = "low";

cyclonev_lcell_comb \F_ctrl_implicit_dst_eretaddr~1 (
	.dataa(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[11] ),
	.datab(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[12] ),
	.datac(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[13] ),
	.datad(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[14] ),
	.datae(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[15] ),
	.dataf(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[16] ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ctrl_implicit_dst_eretaddr~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ctrl_implicit_dst_eretaddr~1 .extended_lut = "off";
defparam \F_ctrl_implicit_dst_eretaddr~1 .lut_mask = 64'h6996966996696996;
defparam \F_ctrl_implicit_dst_eretaddr~1 .shared_arith = "off";

cyclonev_lcell_comb \F_ctrl_implicit_dst_eretaddr~2 (
	.dataa(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[5] ),
	.datab(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[4] ),
	.datac(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[2] ),
	.datad(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[0] ),
	.datae(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[3] ),
	.dataf(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[1] ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ctrl_implicit_dst_eretaddr~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ctrl_implicit_dst_eretaddr~2 .extended_lut = "off";
defparam \F_ctrl_implicit_dst_eretaddr~2 .lut_mask = 64'h9669FFFF6996FFFF;
defparam \F_ctrl_implicit_dst_eretaddr~2 .shared_arith = "off";

cyclonev_lcell_comb \F_ctrl_implicit_dst_eretaddr~0 (
	.dataa(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[5] ),
	.datab(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[4] ),
	.datac(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[2] ),
	.datad(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[1] ),
	.datae(!\F_ctrl_implicit_dst_eretaddr~1_combout ),
	.dataf(!\F_ctrl_implicit_dst_eretaddr~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ctrl_implicit_dst_eretaddr~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ctrl_implicit_dst_eretaddr~0 .extended_lut = "off";
defparam \F_ctrl_implicit_dst_eretaddr~0 .lut_mask = 64'hFFEFFFFFFFFFFFFF;
defparam \F_ctrl_implicit_dst_eretaddr~0 .shared_arith = "off";

dffeas D_ctrl_implicit_dst_eretaddr(
	.clk(clk_clk),
	.d(\F_ctrl_implicit_dst_eretaddr~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_ctrl_implicit_dst_eretaddr~q ),
	.prn(vcc));
defparam D_ctrl_implicit_dst_eretaddr.is_wysiwyg = "true";
defparam D_ctrl_implicit_dst_eretaddr.power_up = "low";

cyclonev_lcell_comb \D_dst_regnum[1]~0 (
	.dataa(!\D_ctrl_b_is_dst~q ),
	.datab(!\D_iw[23]~q ),
	.datac(!\D_iw[18]~q ),
	.datad(!\D_ctrl_implicit_dst_retaddr~q ),
	.datae(!\D_ctrl_implicit_dst_eretaddr~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_dst_regnum[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_dst_regnum[1]~0 .extended_lut = "off";
defparam \D_dst_regnum[1]~0 .lut_mask = 64'hBFFF1FFFBFFF1FFF;
defparam \D_dst_regnum[1]~0 .shared_arith = "off";

dffeas \D_iw[21] (
	.clk(clk_clk),
	.d(\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[21] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_iw[21]~q ),
	.prn(vcc));
defparam \D_iw[21] .is_wysiwyg = "true";
defparam \D_iw[21] .power_up = "low";

cyclonev_lcell_comb \D_dst_regnum[4]~1 (
	.dataa(!\D_ctrl_b_is_dst~q ),
	.datab(!\D_iw[26]~q ),
	.datac(!\D_iw[21]~q ),
	.datad(!\D_ctrl_implicit_dst_retaddr~q ),
	.datae(!\D_ctrl_implicit_dst_eretaddr~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_dst_regnum[4]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_dst_regnum[4]~1 .extended_lut = "off";
defparam \D_dst_regnum[4]~1 .lut_mask = 64'h27FFFFFF27FFFFFF;
defparam \D_dst_regnum[4]~1 .shared_arith = "off";

cyclonev_lcell_comb F_ctrl_ignore_dst(
	.dataa(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[1] ),
	.datab(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[0] ),
	.datac(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[2] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ctrl_ignore_dst~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam F_ctrl_ignore_dst.extended_lut = "off";
defparam F_ctrl_ignore_dst.lut_mask = 64'h6F6F6F6F6F6F6F6F;
defparam F_ctrl_ignore_dst.shared_arith = "off";

dffeas D_ctrl_ignore_dst(
	.clk(clk_clk),
	.d(\F_ctrl_ignore_dst~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_ctrl_ignore_dst~q ),
	.prn(vcc));
defparam D_ctrl_ignore_dst.is_wysiwyg = "true";
defparam D_ctrl_ignore_dst.power_up = "low";

dffeas \D_iw[17] (
	.clk(clk_clk),
	.d(\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[17] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_iw[17]~q ),
	.prn(vcc));
defparam \D_iw[17] .is_wysiwyg = "true";
defparam \D_iw[17] .power_up = "low";

cyclonev_lcell_comb \D_dst_regnum[0]~2 (
	.dataa(!\D_ctrl_b_is_dst~q ),
	.datab(!\D_iw[22]~q ),
	.datac(!\D_iw[17]~q ),
	.datad(!\D_ctrl_implicit_dst_retaddr~q ),
	.datae(!\D_ctrl_implicit_dst_eretaddr~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_dst_regnum[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_dst_regnum[0]~2 .extended_lut = "off";
defparam \D_dst_regnum[0]~2 .lut_mask = 64'h27FFFFFF27FFFFFF;
defparam \D_dst_regnum[0]~2 .shared_arith = "off";

dffeas \D_iw[19] (
	.clk(clk_clk),
	.d(\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[19] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_iw[19]~q ),
	.prn(vcc));
defparam \D_iw[19] .is_wysiwyg = "true";
defparam \D_iw[19] .power_up = "low";

cyclonev_lcell_comb \D_dst_regnum[2]~3 (
	.dataa(!\D_ctrl_b_is_dst~q ),
	.datab(!\D_iw[24]~q ),
	.datac(!\D_iw[19]~q ),
	.datad(!\D_ctrl_implicit_dst_retaddr~q ),
	.datae(!\D_ctrl_implicit_dst_eretaddr~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_dst_regnum[2]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_dst_regnum[2]~3 .extended_lut = "off";
defparam \D_dst_regnum[2]~3 .lut_mask = 64'h27FFFFFF27FFFFFF;
defparam \D_dst_regnum[2]~3 .shared_arith = "off";

dffeas \D_iw[20] (
	.clk(clk_clk),
	.d(\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[20] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_iw[20]~q ),
	.prn(vcc));
defparam \D_iw[20] .is_wysiwyg = "true";
defparam \D_iw[20] .power_up = "low";

cyclonev_lcell_comb \D_dst_regnum[3]~4 (
	.dataa(!\D_ctrl_b_is_dst~q ),
	.datab(!\D_iw[25]~q ),
	.datac(!\D_iw[20]~q ),
	.datad(!\D_ctrl_implicit_dst_retaddr~q ),
	.datae(!\D_ctrl_implicit_dst_eretaddr~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_dst_regnum[3]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_dst_regnum[3]~4 .extended_lut = "off";
defparam \D_dst_regnum[3]~4 .lut_mask = 64'h27FFFFFF27FFFFFF;
defparam \D_dst_regnum[3]~4 .shared_arith = "off";

cyclonev_lcell_comb \Equal302~0 (
	.dataa(!\D_dst_regnum[0]~2_combout ),
	.datab(!\D_dst_regnum[2]~3_combout ),
	.datac(!\D_dst_regnum[3]~4_combout ),
	.datad(!\D_dst_regnum[4]~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal302~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal302~0 .extended_lut = "off";
defparam \Equal302~0 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \Equal302~0 .shared_arith = "off";

cyclonev_lcell_comb D_wr_dst_reg(
	.dataa(!\D_ctrl_ignore_dst~q ),
	.datab(!\D_dst_regnum[1]~0_combout ),
	.datac(!\D_valid~combout ),
	.datad(!\Equal302~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_wr_dst_reg~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam D_wr_dst_reg.extended_lut = "off";
defparam D_wr_dst_reg.lut_mask = 64'hFFBFFFBFFFBFFFBF;
defparam D_wr_dst_reg.shared_arith = "off";

cyclonev_lcell_comb \D_regnum_b_cmp_F~0 (
	.dataa(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[22] ),
	.datab(!\D_dst_regnum[0]~2_combout ),
	.datac(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[24] ),
	.datad(!\D_dst_regnum[2]~3_combout ),
	.datae(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[25] ),
	.dataf(!\D_dst_regnum[3]~4_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_regnum_b_cmp_F~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_regnum_b_cmp_F~0 .extended_lut = "off";
defparam \D_regnum_b_cmp_F~0 .lut_mask = 64'h6996966996696996;
defparam \D_regnum_b_cmp_F~0 .shared_arith = "off";

cyclonev_lcell_comb D_regnum_b_cmp_F(
	.dataa(!\D_dst_regnum[1]~0_combout ),
	.datab(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[23] ),
	.datac(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[26] ),
	.datad(!\D_dst_regnum[4]~1_combout ),
	.datae(!\D_wr_dst_reg~combout ),
	.dataf(!\D_regnum_b_cmp_F~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_regnum_b_cmp_F~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam D_regnum_b_cmp_F.extended_lut = "off";
defparam D_regnum_b_cmp_F.lut_mask = 64'h6996FFFFFFFFFFFF;
defparam D_regnum_b_cmp_F.shared_arith = "off";

dffeas E_regnum_b_cmp_D(
	.clk(clk_clk),
	.d(\D_regnum_b_cmp_F~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\F_stall~0_combout ),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_regnum_b_cmp_D~q ),
	.prn(vcc));
defparam E_regnum_b_cmp_D.is_wysiwyg = "true";
defparam E_regnum_b_cmp_D.power_up = "low";

dffeas A_pipe_flush(
	.clk(clk_clk),
	.d(\A_pipe_flush_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_pipe_flush~q ),
	.prn(vcc));
defparam A_pipe_flush.is_wysiwyg = "true";
defparam A_pipe_flush.power_up = "low";

cyclonev_lcell_comb \Equal149~0 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[13]~q ),
	.datad(!\D_iw[14]~q ),
	.datae(!\D_iw[15]~q ),
	.dataf(!\D_iw[16]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal149~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal149~0 .extended_lut = "off";
defparam \Equal149~0 .lut_mask = 64'hFFFFDFFFFFFFFFFF;
defparam \Equal149~0 .shared_arith = "off";

cyclonev_lcell_comb E_ctrl_trap_inst_nxt(
	.dataa(!\Equal149~0_combout ),
	.datab(!\Equal95~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_ctrl_trap_inst_nxt~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam E_ctrl_trap_inst_nxt.extended_lut = "off";
defparam E_ctrl_trap_inst_nxt.lut_mask = 64'h7777777777777777;
defparam E_ctrl_trap_inst_nxt.shared_arith = "off";

dffeas E_ctrl_trap_inst(
	.clk(clk_clk),
	.d(\E_ctrl_trap_inst_nxt~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_ctrl_trap_inst~q ),
	.prn(vcc));
defparam E_ctrl_trap_inst.is_wysiwyg = "true";
defparam E_ctrl_trap_inst.power_up = "low";

dffeas M_exc_trap_inst_pri15(
	.clk(clk_clk),
	.d(\E_ctrl_trap_inst~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_exc_trap_inst_pri15~q ),
	.prn(vcc));
defparam M_exc_trap_inst_pri15.is_wysiwyg = "true";
defparam M_exc_trap_inst_pri15.power_up = "low";

cyclonev_lcell_comb \D_ctrl_unimp_trap~0 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[14]~q ),
	.datad(!\D_iw[15]~q ),
	.datae(!\D_iw[16]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_unimp_trap~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_unimp_trap~0 .extended_lut = "off";
defparam \D_ctrl_unimp_trap~0 .lut_mask = 64'hFDF7F7FDFDF7F7FD;
defparam \D_ctrl_unimp_trap~0 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_unimp_trap~1 (
	.dataa(!\D_iw[13]~q ),
	.datab(!\Equal95~0_combout ),
	.datac(!\D_ctrl_unimp_trap~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_unimp_trap~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_unimp_trap~1 .extended_lut = "off";
defparam \D_ctrl_unimp_trap~1 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \D_ctrl_unimp_trap~1 .shared_arith = "off";

dffeas E_ctrl_unimp_trap(
	.clk(clk_clk),
	.d(\D_ctrl_unimp_trap~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_ctrl_unimp_trap~q ),
	.prn(vcc));
defparam E_ctrl_unimp_trap.is_wysiwyg = "true";
defparam E_ctrl_unimp_trap.power_up = "low";

dffeas M_exc_unimp_inst_pri15(
	.clk(clk_clk),
	.d(\E_ctrl_unimp_trap~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_exc_unimp_inst_pri15~q ),
	.prn(vcc));
defparam M_exc_unimp_inst_pri15.is_wysiwyg = "true";
defparam M_exc_unimp_inst_pri15.power_up = "low";

dffeas \E_iw[15] (
	.clk(clk_clk),
	.d(\D_iw[15]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_iw[15]~q ),
	.prn(vcc));
defparam \E_iw[15] .is_wysiwyg = "true";
defparam \E_iw[15] .power_up = "low";

dffeas \E_iw[14] (
	.clk(clk_clk),
	.d(\D_iw[14]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_iw[14]~q ),
	.prn(vcc));
defparam \E_iw[14] .is_wysiwyg = "true";
defparam \E_iw[14] .power_up = "low";

dffeas \E_iw[12] (
	.clk(clk_clk),
	.d(\D_iw[12]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_iw[12]~q ),
	.prn(vcc));
defparam \E_iw[12] .is_wysiwyg = "true";
defparam \E_iw[12] .power_up = "low";

dffeas \E_iw[11] (
	.clk(clk_clk),
	.d(\D_iw[11]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_iw[11]~q ),
	.prn(vcc));
defparam \E_iw[11] .is_wysiwyg = "true";
defparam \E_iw[11] .power_up = "low";

dffeas \E_iw[16] (
	.clk(clk_clk),
	.d(\D_iw[16]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_iw[16]~q ),
	.prn(vcc));
defparam \E_iw[16] .is_wysiwyg = "true";
defparam \E_iw[16] .power_up = "low";

dffeas \E_iw[13] (
	.clk(clk_clk),
	.d(\D_iw[13]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_iw[13]~q ),
	.prn(vcc));
defparam \E_iw[13] .is_wysiwyg = "true";
defparam \E_iw[13] .power_up = "low";

dffeas \E_iw[1] (
	.clk(clk_clk),
	.d(\D_iw[1]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_iw[1]~q ),
	.prn(vcc));
defparam \E_iw[1] .is_wysiwyg = "true";
defparam \E_iw[1] .power_up = "low";

dffeas \E_iw[2] (
	.clk(clk_clk),
	.d(\D_iw[2]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_iw[2]~q ),
	.prn(vcc));
defparam \E_iw[2] .is_wysiwyg = "true";
defparam \E_iw[2] .power_up = "low";

dffeas \E_iw[0] (
	.clk(clk_clk),
	.d(\D_iw[0]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_iw[0]~q ),
	.prn(vcc));
defparam \E_iw[0] .is_wysiwyg = "true";
defparam \E_iw[0] .power_up = "low";

dffeas \E_iw[5] (
	.clk(clk_clk),
	.d(\D_iw[5]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_iw[5]~q ),
	.prn(vcc));
defparam \E_iw[5] .is_wysiwyg = "true";
defparam \E_iw[5] .power_up = "low";

dffeas \E_iw[4] (
	.clk(clk_clk),
	.d(\D_iw[4]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_iw[4]~q ),
	.prn(vcc));
defparam \E_iw[4] .is_wysiwyg = "true";
defparam \E_iw[4] .power_up = "low";

dffeas \E_iw[3] (
	.clk(clk_clk),
	.d(\D_iw[3]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_iw[3]~q ),
	.prn(vcc));
defparam \E_iw[3] .is_wysiwyg = "true";
defparam \E_iw[3] .power_up = "low";

cyclonev_lcell_comb \Equal239~0 (
	.dataa(!\E_iw[1]~q ),
	.datab(!\E_iw[2]~q ),
	.datac(!\E_iw[0]~q ),
	.datad(!\E_iw[5]~q ),
	.datae(!\E_iw[4]~q ),
	.dataf(!\E_iw[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal239~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal239~0 .extended_lut = "off";
defparam \Equal239~0 .lut_mask = 64'hFDFFFFFFFFFFFFFF;
defparam \Equal239~0 .shared_arith = "off";

cyclonev_lcell_comb \E_op_rdctl~0 (
	.dataa(!\E_iw[11]~q ),
	.datab(!\E_iw[16]~q ),
	.datac(!\E_iw[13]~q ),
	.datad(!\Equal239~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_op_rdctl~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_op_rdctl~0 .extended_lut = "off";
defparam \E_op_rdctl~0 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \E_op_rdctl~0 .shared_arith = "off";

cyclonev_lcell_comb E_op_break(
	.dataa(!\E_iw[15]~q ),
	.datab(!\E_iw[14]~q ),
	.datac(!\E_iw[12]~q ),
	.datad(!\E_op_rdctl~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_op_break~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam E_op_break.extended_lut = "off";
defparam E_op_break.lut_mask = 64'hFDFFFDFFFDFFFDFF;
defparam E_op_break.shared_arith = "off";

dffeas M_exc_break_inst_pri15(
	.clk(clk_clk),
	.d(\E_op_break~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_exc_break_inst_pri15~q ),
	.prn(vcc));
defparam M_exc_break_inst_pri15.is_wysiwyg = "true";
defparam M_exc_break_inst_pri15.power_up = "low";

cyclonev_lcell_comb \D_ctrl_illegal~0 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[13]~q ),
	.datad(!\D_iw[14]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_illegal~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_illegal~0 .extended_lut = "off";
defparam \D_ctrl_illegal~0 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \D_ctrl_illegal~0 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_illegal~3 (
	.dataa(!\D_iw[16]~q ),
	.datab(!\D_iw[15]~q ),
	.datac(!\D_iw[14]~q ),
	.datad(!\D_iw[13]~q ),
	.datae(!\D_iw[12]~q ),
	.dataf(!\D_iw[11]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_illegal~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_illegal~3 .extended_lut = "off";
defparam \D_ctrl_illegal~3 .lut_mask = 64'h6996966996696996;
defparam \D_ctrl_illegal~3 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_illegal~1 (
	.dataa(!\D_iw[15]~q ),
	.datab(!\D_iw[16]~q ),
	.datac(!\Equal95~0_combout ),
	.datad(!\D_ctrl_illegal~0_combout ),
	.datae(!\D_ctrl_illegal~3_combout ),
	.dataf(!\D_ctrl_flush_pipe_always~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_illegal~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_illegal~1 .extended_lut = "off";
defparam \D_ctrl_illegal~1 .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \D_ctrl_illegal~1 .shared_arith = "off";

dffeas E_ctrl_illegal(
	.clk(clk_clk),
	.d(\D_ctrl_illegal~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_ctrl_illegal~q ),
	.prn(vcc));
defparam E_ctrl_illegal.is_wysiwyg = "true";
defparam E_ctrl_illegal.power_up = "low";

dffeas M_exc_illegal_inst_pri15(
	.clk(clk_clk),
	.d(\E_ctrl_illegal~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_exc_illegal_inst_pri15~q ),
	.prn(vcc));
defparam M_exc_illegal_inst_pri15.is_wysiwyg = "true";
defparam M_exc_illegal_inst_pri15.power_up = "low";

cyclonev_lcell_comb \M_exc_any~0 (
	.dataa(!\M_exc_trap_inst_pri15~q ),
	.datab(!\M_exc_unimp_inst_pri15~q ),
	.datac(!\M_exc_break_inst_pri15~q ),
	.datad(!\M_exc_illegal_inst_pri15~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_exc_any~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_exc_any~0 .extended_lut = "off";
defparam \M_exc_any~0 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \M_exc_any~0 .shared_arith = "off";

dffeas E_wr_dst_reg_from_D(
	.clk(clk_clk),
	.d(\D_wr_dst_reg~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_wr_dst_reg_from_D~q ),
	.prn(vcc));
defparam E_wr_dst_reg_from_D.is_wysiwyg = "true";
defparam E_wr_dst_reg_from_D.power_up = "low";

cyclonev_lcell_comb E_wr_dst_reg(
	.dataa(!\M_pipe_flush~q ),
	.datab(!\E_wr_dst_reg_from_D~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_wr_dst_reg~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam E_wr_dst_reg.extended_lut = "off";
defparam E_wr_dst_reg.lut_mask = 64'h7777777777777777;
defparam E_wr_dst_reg.shared_arith = "off";

dffeas M_wr_dst_reg_from_E(
	.clk(clk_clk),
	.d(\E_wr_dst_reg~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_wr_dst_reg_from_E~q ),
	.prn(vcc));
defparam M_wr_dst_reg_from_E.is_wysiwyg = "true";
defparam M_wr_dst_reg_from_E.power_up = "low";

cyclonev_lcell_comb \M_wr_dst_reg~0 (
	.dataa(!\M_norm_intr_req~q ),
	.datab(!\hbreak_req~0_combout ),
	.datac(!\A_pipe_flush~q ),
	.datad(!\M_exc_any~0_combout ),
	.datae(!\M_wr_dst_reg_from_E~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_wr_dst_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_wr_dst_reg~0 .extended_lut = "off";
defparam \M_wr_dst_reg~0 .lut_mask = 64'hFFFFFF7FFFFFFF7F;
defparam \M_wr_dst_reg~0 .shared_arith = "off";

dffeas A_wr_dst_reg_from_M(
	.clk(clk_clk),
	.d(\M_wr_dst_reg~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_wr_dst_reg_from_M~q ),
	.prn(vcc));
defparam A_wr_dst_reg_from_M.is_wysiwyg = "true";
defparam A_wr_dst_reg_from_M.power_up = "low";

cyclonev_lcell_comb \A_wr_dst_reg~0 (
	.dataa(!\A_exc_any~q ),
	.datab(!\A_exc_allowed~q ),
	.datac(!\A_wr_dst_reg_from_M~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_dst_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_dst_reg~0 .extended_lut = "off";
defparam \A_wr_dst_reg~0 .lut_mask = 64'hF7F7F7F7F7F7F7F7;
defparam \A_wr_dst_reg~0 .shared_arith = "off";

cyclonev_lcell_comb \M_exc_break~0 (
	.dataa(!\M_exc_break_inst_pri15~q ),
	.datab(!\M_norm_intr_req~q ),
	.datac(!\hbreak_req~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_exc_break~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_exc_break~0 .extended_lut = "off";
defparam \M_exc_break~0 .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \M_exc_break~0 .shared_arith = "off";

dffeas A_exc_break(
	.clk(clk_clk),
	.d(\M_exc_break~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_exc_break~q ),
	.prn(vcc));
defparam A_exc_break.is_wysiwyg = "true";
defparam A_exc_break.power_up = "low";

dffeas \E_dst_regnum[0] (
	.clk(clk_clk),
	.d(\D_dst_regnum[0]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_dst_regnum[0]~q ),
	.prn(vcc));
defparam \E_dst_regnum[0] .is_wysiwyg = "true";
defparam \E_dst_regnum[0] .power_up = "low";

dffeas \M_dst_regnum[0] (
	.clk(clk_clk),
	.d(\E_dst_regnum[0]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_dst_regnum[0]~q ),
	.prn(vcc));
defparam \M_dst_regnum[0] .is_wysiwyg = "true";
defparam \M_dst_regnum[0] .power_up = "low";

dffeas \A_dst_regnum_from_M[0] (
	.clk(clk_clk),
	.d(\M_dst_regnum[0]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_dst_regnum_from_M[0]~q ),
	.prn(vcc));
defparam \A_dst_regnum_from_M[0] .is_wysiwyg = "true";
defparam \A_dst_regnum_from_M[0] .power_up = "low";

cyclonev_lcell_comb \A_dst_regnum~0 (
	.dataa(!\A_exc_any~q ),
	.datab(!\A_exc_break~q ),
	.datac(!\A_dst_regnum_from_M[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dst_regnum~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dst_regnum~0 .extended_lut = "off";
defparam \A_dst_regnum~0 .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \A_dst_regnum~0 .shared_arith = "off";

dffeas \E_dst_regnum[1] (
	.clk(clk_clk),
	.d(\D_dst_regnum[1]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_dst_regnum[1]~q ),
	.prn(vcc));
defparam \E_dst_regnum[1] .is_wysiwyg = "true";
defparam \E_dst_regnum[1] .power_up = "low";

dffeas \M_dst_regnum[1] (
	.clk(clk_clk),
	.d(\E_dst_regnum[1]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_dst_regnum[1]~q ),
	.prn(vcc));
defparam \M_dst_regnum[1] .is_wysiwyg = "true";
defparam \M_dst_regnum[1] .power_up = "low";

dffeas \A_dst_regnum_from_M[1] (
	.clk(clk_clk),
	.d(\M_dst_regnum[1]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_dst_regnum_from_M[1]~q ),
	.prn(vcc));
defparam \A_dst_regnum_from_M[1] .is_wysiwyg = "true";
defparam \A_dst_regnum_from_M[1] .power_up = "low";

cyclonev_lcell_comb \A_dst_regnum~1 (
	.dataa(!\A_exc_any~q ),
	.datab(!\A_exc_break~q ),
	.datac(!\A_dst_regnum_from_M[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dst_regnum~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dst_regnum~1 .extended_lut = "off";
defparam \A_dst_regnum~1 .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \A_dst_regnum~1 .shared_arith = "off";

dffeas \E_dst_regnum[2] (
	.clk(clk_clk),
	.d(\D_dst_regnum[2]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_dst_regnum[2]~q ),
	.prn(vcc));
defparam \E_dst_regnum[2] .is_wysiwyg = "true";
defparam \E_dst_regnum[2] .power_up = "low";

dffeas \M_dst_regnum[2] (
	.clk(clk_clk),
	.d(\E_dst_regnum[2]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_dst_regnum[2]~q ),
	.prn(vcc));
defparam \M_dst_regnum[2] .is_wysiwyg = "true";
defparam \M_dst_regnum[2] .power_up = "low";

dffeas \A_dst_regnum_from_M[2] (
	.clk(clk_clk),
	.d(\M_dst_regnum[2]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_dst_regnum_from_M[2]~q ),
	.prn(vcc));
defparam \A_dst_regnum_from_M[2] .is_wysiwyg = "true";
defparam \A_dst_regnum_from_M[2] .power_up = "low";

cyclonev_lcell_comb \A_dst_regnum~2 (
	.dataa(!\A_exc_any~q ),
	.datab(!\A_exc_break~q ),
	.datac(!\A_dst_regnum_from_M[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dst_regnum~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dst_regnum~2 .extended_lut = "off";
defparam \A_dst_regnum~2 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \A_dst_regnum~2 .shared_arith = "off";

cyclonev_lcell_comb \A_regnum_b_cmp_F~0 (
	.dataa(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[23] ),
	.datab(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[24] ),
	.datac(!\A_dst_regnum~1_combout ),
	.datad(!\A_dst_regnum~2_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_regnum_b_cmp_F~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_regnum_b_cmp_F~0 .extended_lut = "off";
defparam \A_regnum_b_cmp_F~0 .lut_mask = 64'h6996699669966996;
defparam \A_regnum_b_cmp_F~0 .shared_arith = "off";

dffeas \E_dst_regnum[3] (
	.clk(clk_clk),
	.d(\D_dst_regnum[3]~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_dst_regnum[3]~q ),
	.prn(vcc));
defparam \E_dst_regnum[3] .is_wysiwyg = "true";
defparam \E_dst_regnum[3] .power_up = "low";

dffeas \M_dst_regnum[3] (
	.clk(clk_clk),
	.d(\E_dst_regnum[3]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_dst_regnum[3]~q ),
	.prn(vcc));
defparam \M_dst_regnum[3] .is_wysiwyg = "true";
defparam \M_dst_regnum[3] .power_up = "low";

dffeas \A_dst_regnum_from_M[3] (
	.clk(clk_clk),
	.d(\M_dst_regnum[3]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_dst_regnum_from_M[3]~q ),
	.prn(vcc));
defparam \A_dst_regnum_from_M[3] .is_wysiwyg = "true";
defparam \A_dst_regnum_from_M[3] .power_up = "low";

cyclonev_lcell_comb \A_dst_regnum~3 (
	.dataa(!\A_exc_any~q ),
	.datab(!\A_exc_break~q ),
	.datac(!\A_dst_regnum_from_M[3]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dst_regnum~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dst_regnum~3 .extended_lut = "off";
defparam \A_dst_regnum~3 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \A_dst_regnum~3 .shared_arith = "off";

dffeas \E_dst_regnum[4] (
	.clk(clk_clk),
	.d(\D_dst_regnum[4]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_dst_regnum[4]~q ),
	.prn(vcc));
defparam \E_dst_regnum[4] .is_wysiwyg = "true";
defparam \E_dst_regnum[4] .power_up = "low";

dffeas \M_dst_regnum[4] (
	.clk(clk_clk),
	.d(\E_dst_regnum[4]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_dst_regnum[4]~q ),
	.prn(vcc));
defparam \M_dst_regnum[4] .is_wysiwyg = "true";
defparam \M_dst_regnum[4] .power_up = "low";

dffeas \A_dst_regnum_from_M[4] (
	.clk(clk_clk),
	.d(\M_dst_regnum[4]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_dst_regnum_from_M[4]~q ),
	.prn(vcc));
defparam \A_dst_regnum_from_M[4] .is_wysiwyg = "true";
defparam \A_dst_regnum_from_M[4] .power_up = "low";

cyclonev_lcell_comb \A_dst_regnum~4 (
	.dataa(!\A_exc_any~q ),
	.datab(!\A_exc_break~q ),
	.datac(!\A_dst_regnum_from_M[4]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dst_regnum~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dst_regnum~4 .extended_lut = "off";
defparam \A_dst_regnum~4 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \A_dst_regnum~4 .shared_arith = "off";

cyclonev_lcell_comb \A_regnum_b_cmp_F~1 (
	.dataa(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[25] ),
	.datab(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[26] ),
	.datac(!\A_dst_regnum~3_combout ),
	.datad(!\A_dst_regnum~4_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_regnum_b_cmp_F~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_regnum_b_cmp_F~1 .extended_lut = "off";
defparam \A_regnum_b_cmp_F~1 .lut_mask = 64'h6996699669966996;
defparam \A_regnum_b_cmp_F~1 .shared_arith = "off";

cyclonev_lcell_comb A_regnum_b_cmp_F(
	.dataa(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[22] ),
	.datab(!\A_wr_dst_reg~0_combout ),
	.datac(!\A_dst_regnum~0_combout ),
	.datad(!\A_regnum_b_cmp_F~0_combout ),
	.datae(!\A_regnum_b_cmp_F~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_regnum_b_cmp_F~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam A_regnum_b_cmp_F.extended_lut = "off";
defparam A_regnum_b_cmp_F.lut_mask = 64'h7BFFFFFF7BFFFFFF;
defparam A_regnum_b_cmp_F.shared_arith = "off";

cyclonev_lcell_comb \M_regnum_b_cmp_F~0 (
	.dataa(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[22] ),
	.datab(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[23] ),
	.datac(!\M_dst_regnum[0]~q ),
	.datad(!\M_dst_regnum[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_regnum_b_cmp_F~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_regnum_b_cmp_F~0 .extended_lut = "off";
defparam \M_regnum_b_cmp_F~0 .lut_mask = 64'h6996699669966996;
defparam \M_regnum_b_cmp_F~0 .shared_arith = "off";

cyclonev_lcell_comb \M_regnum_b_cmp_F~1 (
	.dataa(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[25] ),
	.datab(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[26] ),
	.datac(!\M_dst_regnum[3]~q ),
	.datad(!\M_dst_regnum[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_regnum_b_cmp_F~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_regnum_b_cmp_F~1 .extended_lut = "off";
defparam \M_regnum_b_cmp_F~1 .lut_mask = 64'h6996699669966996;
defparam \M_regnum_b_cmp_F~1 .shared_arith = "off";

cyclonev_lcell_comb M_regnum_b_cmp_F(
	.dataa(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[24] ),
	.datab(!\M_dst_regnum[2]~q ),
	.datac(!\M_wr_dst_reg~0_combout ),
	.datad(!\M_regnum_b_cmp_F~0_combout ),
	.datae(!\M_regnum_b_cmp_F~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_regnum_b_cmp_F~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam M_regnum_b_cmp_F.extended_lut = "off";
defparam M_regnum_b_cmp_F.lut_mask = 64'hF6FFFFFFF6FFFFFF;
defparam M_regnum_b_cmp_F.shared_arith = "off";

cyclonev_lcell_comb \E_regnum_b_cmp_F~0 (
	.dataa(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[22] ),
	.datab(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[23] ),
	.datac(!\E_wr_dst_reg~combout ),
	.datad(!\E_dst_regnum[0]~q ),
	.datae(!\E_dst_regnum[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_regnum_b_cmp_F~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_regnum_b_cmp_F~0 .extended_lut = "off";
defparam \E_regnum_b_cmp_F~0 .lut_mask = 64'h6F9F9F6F6F9F9F6F;
defparam \E_regnum_b_cmp_F~0 .shared_arith = "off";

cyclonev_lcell_comb \E_regnum_b_cmp_F~1 (
	.dataa(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[24] ),
	.datab(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[25] ),
	.datac(!\E_dst_regnum[2]~q ),
	.datad(!\E_dst_regnum[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_regnum_b_cmp_F~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_regnum_b_cmp_F~1 .extended_lut = "off";
defparam \E_regnum_b_cmp_F~1 .lut_mask = 64'h6996699669966996;
defparam \E_regnum_b_cmp_F~1 .shared_arith = "off";

cyclonev_lcell_comb E_regnum_b_cmp_F(
	.dataa(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[26] ),
	.datab(!\E_dst_regnum[4]~q ),
	.datac(!\E_regnum_b_cmp_F~0_combout ),
	.datad(!\E_regnum_b_cmp_F~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_regnum_b_cmp_F~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam E_regnum_b_cmp_F.extended_lut = "off";
defparam E_regnum_b_cmp_F.lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam E_regnum_b_cmp_F.shared_arith = "off";

dffeas M_regnum_b_cmp_D(
	.clk(clk_clk),
	.d(\E_regnum_b_cmp_F~combout ),
	.asdata(\E_regnum_b_cmp_D~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\F_stall~0_combout ),
	.ena(!\A_mem_stall~q ),
	.q(\M_regnum_b_cmp_D~q ),
	.prn(vcc));
defparam M_regnum_b_cmp_D.is_wysiwyg = "true";
defparam M_regnum_b_cmp_D.power_up = "low";

dffeas A_regnum_b_cmp_D(
	.clk(clk_clk),
	.d(\M_regnum_b_cmp_F~combout ),
	.asdata(\M_regnum_b_cmp_D~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\F_stall~0_combout ),
	.ena(!\A_mem_stall~q ),
	.q(\A_regnum_b_cmp_D~q ),
	.prn(vcc));
defparam A_regnum_b_cmp_D.is_wysiwyg = "true";
defparam A_regnum_b_cmp_D.power_up = "low";

dffeas W_regnum_b_cmp_D(
	.clk(clk_clk),
	.d(\A_regnum_b_cmp_F~combout ),
	.asdata(\A_regnum_b_cmp_D~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\F_stall~0_combout ),
	.ena(vcc),
	.q(\W_regnum_b_cmp_D~q ),
	.prn(vcc));
defparam W_regnum_b_cmp_D.is_wysiwyg = "true";
defparam W_regnum_b_cmp_D.power_up = "low";

cyclonev_lcell_comb \D_src2_reg[0]~0 (
	.dataa(!\D_ctrl_b_is_dst~q ),
	.datab(!\E_regnum_b_cmp_D~q ),
	.datac(!\W_regnum_b_cmp_D~q ),
	.datad(!\A_regnum_b_cmp_D~q ),
	.datae(!\M_regnum_b_cmp_D~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[0]~0 .extended_lut = "off";
defparam \D_src2_reg[0]~0 .lut_mask = 64'hEFFFFFFFEFFFFFFF;
defparam \D_src2_reg[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[0]~4 (
	.dataa(!\Equal304~0_combout ),
	.datab(!\D_src2_reg[0]~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[0]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[0]~4 .extended_lut = "off";
defparam \D_src2_reg[0]~4 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \D_src2_reg[0]~4 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[0]~1 (
	.dataa(!\D_ctrl_b_is_dst~q ),
	.datab(!\E_regnum_b_cmp_D~q ),
	.datac(!\W_regnum_b_cmp_D~q ),
	.datad(!\A_regnum_b_cmp_D~q ),
	.datae(!\M_regnum_b_cmp_D~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[0]~1 .extended_lut = "off";
defparam \D_src2_reg[0]~1 .lut_mask = 64'hBFFFFFFFBFFFFFFF;
defparam \D_src2_reg[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[0]~5 (
	.dataa(!\Equal304~0_combout ),
	.datab(!\D_src2_reg[0]~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[0]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[0]~5 .extended_lut = "off";
defparam \D_src2_reg[0]~5 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \D_src2_reg[0]~5 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[0]~6 (
	.dataa(!\D_src2_reg[0]~4_combout ),
	.datab(!\D_src2_reg[0]~5_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[0]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[0]~6 .extended_lut = "off";
defparam \D_src2_reg[0]~6 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \D_src2_reg[0]~6 .shared_arith = "off";

cyclonev_lcell_comb \F_ctrl_src2_choose_imm~1 (
	.dataa(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[13] ),
	.datab(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[4] ),
	.datac(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[3] ),
	.datad(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[2] ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ctrl_src2_choose_imm~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ctrl_src2_choose_imm~1 .extended_lut = "off";
defparam \F_ctrl_src2_choose_imm~1 .lut_mask = 64'hFFBFFFBFFFBFFFBF;
defparam \F_ctrl_src2_choose_imm~1 .shared_arith = "off";

cyclonev_lcell_comb \F_ctrl_src2_choose_imm~0 (
	.dataa(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[11] ),
	.datab(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[12] ),
	.datac(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[1] ),
	.datad(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[0] ),
	.datae(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[5] ),
	.dataf(!\F_ctrl_src2_choose_imm~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ctrl_src2_choose_imm~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ctrl_src2_choose_imm~0 .extended_lut = "off";
defparam \F_ctrl_src2_choose_imm~0 .lut_mask = 64'hFBFFFFFFFFFFFFFF;
defparam \F_ctrl_src2_choose_imm~0 .shared_arith = "off";

dffeas D_ctrl_src2_choose_imm(
	.clk(clk_clk),
	.d(\F_ctrl_src2_choose_imm~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_ctrl_src2_choose_imm~q ),
	.prn(vcc));
defparam D_ctrl_src2_choose_imm.is_wysiwyg = "true";
defparam D_ctrl_src2_choose_imm.power_up = "low";

cyclonev_lcell_comb \D_ctrl_logic~0 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[13]~q ),
	.datad(!\D_iw[16]~q ),
	.datae(!\Equal95~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_logic~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_logic~0 .extended_lut = "off";
defparam \D_ctrl_logic~0 .lut_mask = 64'hFFBFFFFFFFBFFFFF;
defparam \D_ctrl_logic~0 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_logic~1 (
	.dataa(!\D_ctrl_logic~0_combout ),
	.datab(!\D_iw[4]~q ),
	.datac(!\D_iw[3]~q ),
	.datad(!\D_iw[2]~q ),
	.datae(!\D_iw[1]~q ),
	.dataf(!\D_iw[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_logic~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_logic~1 .extended_lut = "off";
defparam \D_ctrl_logic~1 .lut_mask = 64'hFFFFFFFFFFFF7FFF;
defparam \D_ctrl_logic~1 .shared_arith = "off";

dffeas E_ctrl_logic(
	.clk(clk_clk),
	.d(\D_ctrl_logic~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_ctrl_logic~q ),
	.prn(vcc));
defparam E_ctrl_logic.is_wysiwyg = "true";
defparam E_ctrl_logic.power_up = "low";

cyclonev_lcell_comb \Equal95~4 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[1]~q ),
	.datac(!\D_iw[2]~q ),
	.datad(!\D_iw[3]~q ),
	.datae(!\D_iw[4]~q ),
	.dataf(!\D_iw[5]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal95~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal95~4 .extended_lut = "off";
defparam \Equal95~4 .lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam \Equal95~4 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_retaddr~1 (
	.dataa(!\D_iw[16]~q ),
	.datab(!\D_iw[15]~q ),
	.datac(!\D_iw[14]~q ),
	.datad(!\D_iw[13]~q ),
	.datae(!\D_iw[12]~q ),
	.dataf(!\D_iw[11]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_retaddr~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_retaddr~1 .extended_lut = "off";
defparam \D_ctrl_retaddr~1 .lut_mask = 64'h7BFFB7FFB7FF7BFF;
defparam \D_ctrl_retaddr~1 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_retaddr~0 (
	.dataa(!\Equal149~0_combout ),
	.datab(!\Equal95~0_combout ),
	.datac(!\D_ctrl_illegal~3_combout ),
	.datad(!\D_ctrl_flush_pipe_always~2_combout ),
	.datae(!\Equal95~4_combout ),
	.dataf(!\D_ctrl_retaddr~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_retaddr~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_retaddr~0 .extended_lut = "off";
defparam \D_ctrl_retaddr~0 .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \D_ctrl_retaddr~0 .shared_arith = "off";

dffeas E_ctrl_retaddr(
	.clk(clk_clk),
	.d(\D_ctrl_retaddr~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_ctrl_retaddr~q ),
	.prn(vcc));
defparam E_ctrl_retaddr.is_wysiwyg = "true";
defparam E_ctrl_retaddr.power_up = "low";

cyclonev_lcell_comb \E_alu_result~0 (
	.dataa(!\E_ctrl_cmp~q ),
	.datab(!\E_ctrl_logic~q ),
	.datac(!\E_ctrl_retaddr~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result~0 .extended_lut = "off";
defparam \E_alu_result~0 .lut_mask = 64'hFEFEFEFEFEFEFEFE;
defparam \E_alu_result~0 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[0]~2 (
	.dataa(!\Equal304~0_combout ),
	.datab(!\D_src2_reg[0]~0_combout ),
	.datac(!\D_src2_reg[0]~1_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[0]~2 .extended_lut = "off";
defparam \D_src2_reg[0]~2 .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \D_src2_reg[0]~2 .shared_arith = "off";

cyclonev_lcell_comb \D_logic_op_raw[1]~1 (
	.dataa(!\D_iw[15]~q ),
	.datab(!\D_iw[4]~q ),
	.datac(!\Equal95~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_logic_op_raw[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_logic_op_raw[1]~1 .extended_lut = "off";
defparam \D_logic_op_raw[1]~1 .lut_mask = 64'h5353535353535353;
defparam \D_logic_op_raw[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_alu_force_xor~1 (
	.dataa(!\D_iw[5]~q ),
	.datab(!\D_iw[4]~q ),
	.datac(!\D_iw[3]~q ),
	.datad(!\D_iw[2]~q ),
	.datae(!\D_iw[1]~q ),
	.dataf(!\D_iw[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_alu_force_xor~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_alu_force_xor~1 .extended_lut = "off";
defparam \D_ctrl_alu_force_xor~1 .lut_mask = 64'hFFFFFFFFEFDFDFEF;
defparam \D_ctrl_alu_force_xor~1 .shared_arith = "off";

cyclonev_lcell_comb \Equal149~5 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[13]~q ),
	.datad(!\D_iw[14]~q ),
	.datae(!\D_iw[15]~q ),
	.dataf(!\D_iw[16]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal149~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal149~5 .extended_lut = "off";
defparam \Equal149~5 .lut_mask = 64'hFFFFFEFFFFFFFFFF;
defparam \Equal149~5 .shared_arith = "off";

cyclonev_lcell_comb \Equal149~1 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[13]~q ),
	.datad(!\D_iw[14]~q ),
	.datae(!\D_iw[15]~q ),
	.dataf(!\D_iw[16]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal149~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal149~1 .extended_lut = "off";
defparam \Equal149~1 .lut_mask = 64'hFFFFFFFFFEFFFFFF;
defparam \Equal149~1 .shared_arith = "off";

cyclonev_lcell_comb \Equal149~2 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[13]~q ),
	.datad(!\D_iw[14]~q ),
	.datae(!\D_iw[15]~q ),
	.dataf(!\D_iw[16]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal149~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal149~2 .extended_lut = "off";
defparam \Equal149~2 .lut_mask = 64'hFFFFFFFEFFFFFFFF;
defparam \Equal149~2 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_alu_force_xor~0 (
	.dataa(!\Equal95~0_combout ),
	.datab(!\Equal149~4_combout ),
	.datac(!\Equal149~5_combout ),
	.datad(!\Equal149~1_combout ),
	.datae(!\Equal149~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_alu_force_xor~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_alu_force_xor~0 .extended_lut = "off";
defparam \D_ctrl_alu_force_xor~0 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \D_ctrl_alu_force_xor~0 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_alu_force_xor~2 (
	.dataa(!\D_ctrl_alu_force_xor~1_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\D_ctrl_alu_force_xor~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_alu_force_xor~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_alu_force_xor~2 .extended_lut = "off";
defparam \D_ctrl_alu_force_xor~2 .lut_mask = 64'hFFAAFFAAFFAAFFAA;
defparam \D_ctrl_alu_force_xor~2 .shared_arith = "off";

cyclonev_lcell_comb \D_logic_op[1]~0 (
	.dataa(!\D_logic_op_raw[1]~1_combout ),
	.datab(!\D_ctrl_alu_force_xor~2_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_logic_op[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_logic_op[1]~0 .extended_lut = "off";
defparam \D_logic_op[1]~0 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \D_logic_op[1]~0 .shared_arith = "off";

dffeas \E_logic_op[1] (
	.clk(clk_clk),
	.d(\D_logic_op[1]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_logic_op[1]~q ),
	.prn(vcc));
defparam \E_logic_op[1] .is_wysiwyg = "true";
defparam \E_logic_op[1] .power_up = "low";

cyclonev_lcell_comb \D_logic_op_raw[0]~0 (
	.dataa(!\D_iw[14]~q ),
	.datab(!\D_iw[3]~q ),
	.datac(!\Equal95~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_logic_op_raw[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_logic_op_raw[0]~0 .extended_lut = "off";
defparam \D_logic_op_raw[0]~0 .lut_mask = 64'h5353535353535353;
defparam \D_logic_op_raw[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \D_logic_op[0]~1 (
	.dataa(!\D_logic_op_raw[0]~0_combout ),
	.datab(!\D_ctrl_alu_force_xor~2_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_logic_op[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_logic_op[0]~1 .extended_lut = "off";
defparam \D_logic_op[0]~1 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \D_logic_op[0]~1 .shared_arith = "off";

dffeas \E_logic_op[0] (
	.clk(clk_clk),
	.d(\D_logic_op[0]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_logic_op[0]~q ),
	.prn(vcc));
defparam \E_logic_op[0] .is_wysiwyg = "true";
defparam \E_logic_op[0] .power_up = "low";

cyclonev_lcell_comb \E_alu_result~10 (
	.dataa(!\E_src2[31]~q ),
	.datab(!\E_src1[31]~q ),
	.datac(!\E_logic_op[1]~q ),
	.datad(!\E_logic_op[0]~q ),
	.datae(!\E_ctrl_logic~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result~10 .extended_lut = "off";
defparam \E_alu_result~10 .lut_mask = 64'h6996FFFF6996FFFF;
defparam \E_alu_result~10 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[31] (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\Add9~73_sumout ),
	.datac(!\E_alu_result~10_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[31]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[31] .extended_lut = "off";
defparam \E_alu_result[31] .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \E_alu_result[31] .shared_arith = "off";

dffeas \M_alu_result[31] (
	.clk(clk_clk),
	.d(\E_alu_result[31]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_alu_result[31]~q ),
	.prn(vcc));
defparam \M_alu_result[31] .is_wysiwyg = "true";
defparam \M_alu_result[31] .power_up = "low";

cyclonev_lcell_comb \Equal219~0 (
	.dataa(!\E_iw[1]~q ),
	.datab(!\E_iw[2]~q ),
	.datac(!\E_iw[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal219~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal219~0 .extended_lut = "off";
defparam \Equal219~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \Equal219~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal219~1 (
	.dataa(!\E_iw[4]~q ),
	.datab(!\Equal219~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal219~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal219~1 .extended_lut = "off";
defparam \Equal219~1 .lut_mask = 64'h7777777777777777;
defparam \Equal219~1 .shared_arith = "off";

dffeas M_ctrl_ld32(
	.clk(clk_clk),
	.d(\Equal219~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_ctrl_ld32~q ),
	.prn(vcc));
defparam M_ctrl_ld32.is_wysiwyg = "true";
defparam M_ctrl_ld32.power_up = "low";

dffeas A_ctrl_ld32(
	.clk(clk_clk),
	.d(\M_ctrl_ld32~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_ctrl_ld32~q ),
	.prn(vcc));
defparam A_ctrl_ld32.is_wysiwyg = "true";
defparam A_ctrl_ld32.power_up = "low";

dffeas \d_readdata_d1[31] (
	.clk(clk_clk),
	.d(d_readdata[31]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[31]~q ),
	.prn(vcc));
defparam \d_readdata_d1[31] .is_wysiwyg = "true";
defparam \d_readdata_d1[31] .power_up = "low";

dffeas \M_alu_result[1] (
	.clk(clk_clk),
	.d(\E_alu_result[1]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_alu_result[1]~q ),
	.prn(vcc));
defparam \M_alu_result[1] .is_wysiwyg = "true";
defparam \M_alu_result[1] .power_up = "low";

dffeas \d_readdata_d1[1] (
	.clk(clk_clk),
	.d(d_readdata[1]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[1]~q ),
	.prn(vcc));
defparam \d_readdata_d1[1] .is_wysiwyg = "true";
defparam \d_readdata_d1[1] .power_up = "low";

dffeas \d_readdata_d1[17] (
	.clk(clk_clk),
	.d(d_readdata[17]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[17]~q ),
	.prn(vcc));
defparam \d_readdata_d1[17] .is_wysiwyg = "true";
defparam \d_readdata_d1[17] .power_up = "low";

dffeas \d_readdata_d1[9] (
	.clk(clk_clk),
	.d(d_readdata[9]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[9]~q ),
	.prn(vcc));
defparam \d_readdata_d1[9] .is_wysiwyg = "true";
defparam \d_readdata_d1[9] .power_up = "low";

dffeas \d_readdata_d1[25] (
	.clk(clk_clk),
	.d(d_readdata[25]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[25]~q ),
	.prn(vcc));
defparam \d_readdata_d1[25] .is_wysiwyg = "true";
defparam \d_readdata_d1[25] .power_up = "low";

cyclonev_lcell_comb \Equal212~0 (
	.dataa(!\E_iw[1]~q ),
	.datab(!\E_iw[0]~q ),
	.datac(!\E_iw[4]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal212~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal212~0 .extended_lut = "off";
defparam \Equal212~0 .lut_mask = 64'hF7F7F7F7F7F7F7F7;
defparam \Equal212~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal212~1 (
	.dataa(!\E_iw[3]~q ),
	.datab(!\Equal212~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal212~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal212~1 .extended_lut = "off";
defparam \Equal212~1 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \Equal212~1 .shared_arith = "off";

dffeas M_ctrl_ld8(
	.clk(clk_clk),
	.d(\Equal212~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_ctrl_ld8~q ),
	.prn(vcc));
defparam M_ctrl_ld8.is_wysiwyg = "true";
defparam M_ctrl_ld8.power_up = "low";

cyclonev_lcell_comb \Equal215~0 (
	.dataa(!\E_iw[3]~q ),
	.datab(!\Equal212~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal215~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal215~0 .extended_lut = "off";
defparam \Equal215~0 .lut_mask = 64'h7777777777777777;
defparam \Equal215~0 .shared_arith = "off";

dffeas M_ctrl_ld16(
	.clk(clk_clk),
	.d(\Equal215~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_ctrl_ld16~q ),
	.prn(vcc));
defparam M_ctrl_ld16.is_wysiwyg = "true";
defparam M_ctrl_ld16.power_up = "low";

cyclonev_lcell_comb \M_ld_align_sh16~0 (
	.dataa(!\M_exc_any~combout ),
	.datab(!\M_mem_baddr[1]~q ),
	.datac(!\M_ctrl_ld8~q ),
	.datad(!\M_ctrl_ld16~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_ld_align_sh16~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_ld_align_sh16~0 .extended_lut = "off";
defparam \M_ld_align_sh16~0 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \M_ld_align_sh16~0 .shared_arith = "off";

dffeas A_ld_align_sh16(
	.clk(clk_clk),
	.d(\M_ld_align_sh16~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_ld_align_sh16~q ),
	.prn(vcc));
defparam A_ld_align_sh16.is_wysiwyg = "true";
defparam A_ld_align_sh16.power_up = "low";

cyclonev_lcell_comb \F_ctrl_hi_imm16~0 (
	.dataa(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[1] ),
	.datab(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[0] ),
	.datac(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[5] ),
	.datad(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[4] ),
	.datae(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[3] ),
	.dataf(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[2] ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ctrl_hi_imm16~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ctrl_hi_imm16~0 .extended_lut = "off";
defparam \F_ctrl_hi_imm16~0 .lut_mask = 64'hEFFFFFFFFFFFFFFF;
defparam \F_ctrl_hi_imm16~0 .shared_arith = "off";

dffeas D_ctrl_hi_imm16(
	.clk(clk_clk),
	.d(\F_ctrl_hi_imm16~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_ctrl_hi_imm16~q ),
	.prn(vcc));
defparam D_ctrl_hi_imm16.is_wysiwyg = "true";
defparam D_ctrl_hi_imm16.power_up = "low";

cyclonev_lcell_comb \D_ctrl_shift_right_arith~0 (
	.dataa(!\D_iw[12]~q ),
	.datab(!\D_iw[13]~q ),
	.datac(!\Equal95~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_shift_right_arith~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_shift_right_arith~0 .extended_lut = "off";
defparam \D_ctrl_shift_right_arith~0 .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \D_ctrl_shift_right_arith~0 .shared_arith = "off";

cyclonev_lcell_comb \E_src2[1]~0 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\D_ctrl_src2_choose_imm~q ),
	.datac(!\D_ctrl_hi_imm16~q ),
	.datad(!\D_ctrl_shift_right_arith~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_src2[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_src2[1]~0 .extended_lut = "off";
defparam \E_src2[1]~0 .lut_mask = 64'hFF7FFF7FFF7FFF7F;
defparam \E_src2[1]~0 .shared_arith = "off";

dffeas \D_iw[6] (
	.clk(clk_clk),
	.d(\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[6] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_iw[6]~q ),
	.prn(vcc));
defparam \D_iw[6] .is_wysiwyg = "true";
defparam \D_iw[6] .power_up = "low";

dffeas \d_readdata_d1[0] (
	.clk(clk_clk),
	.d(d_readdata[0]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[0]~q ),
	.prn(vcc));
defparam \d_readdata_d1[0] .is_wysiwyg = "true";
defparam \d_readdata_d1[0] .power_up = "low";

dffeas \d_readdata_d1[16] (
	.clk(clk_clk),
	.d(d_readdata[16]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[16]~q ),
	.prn(vcc));
defparam \d_readdata_d1[16] .is_wysiwyg = "true";
defparam \d_readdata_d1[16] .power_up = "low";

dffeas \d_readdata_d1[8] (
	.clk(clk_clk),
	.d(d_readdata[8]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[8]~q ),
	.prn(vcc));
defparam \d_readdata_d1[8] .is_wysiwyg = "true";
defparam \d_readdata_d1[8] .power_up = "low";

dffeas \d_readdata_d1[24] (
	.clk(clk_clk),
	.d(d_readdata[24]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[24]~q ),
	.prn(vcc));
defparam \d_readdata_d1[24] .is_wysiwyg = "true";
defparam \d_readdata_d1[24] .power_up = "low";

cyclonev_lcell_comb \A_slow_inst_result_nxt[0]~0 (
	.dataa(!\d_readdata_d1[0]~q ),
	.datab(!\d_readdata_d1[16]~q ),
	.datac(!\d_readdata_d1[8]~q ),
	.datad(!\d_readdata_d1[24]~q ),
	.datae(!\A_ld_align_sh16~q ),
	.dataf(!\A_ld_align_sh8~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[0]~0 .extended_lut = "off";
defparam \A_slow_inst_result_nxt[0]~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_slow_inst_result_nxt[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_ld~0 (
	.dataa(!\D_iw[4]~q ),
	.datab(!\D_iw[0]~q ),
	.datac(!\D_iw[1]~q ),
	.datad(!\D_iw[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_ld~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_ld~0 .extended_lut = "off";
defparam \D_ctrl_ld~0 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \D_ctrl_ld~0 .shared_arith = "off";

dffeas E_ctrl_ld(
	.clk(clk_clk),
	.d(\D_ctrl_ld~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_ctrl_ld~q ),
	.prn(vcc));
defparam E_ctrl_ld.is_wysiwyg = "true";
defparam E_ctrl_ld.power_up = "low";

dffeas M_ctrl_ld(
	.clk(clk_clk),
	.d(\E_ctrl_ld~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_ctrl_ld~q ),
	.prn(vcc));
defparam M_ctrl_ld.is_wysiwyg = "true";
defparam M_ctrl_ld.power_up = "low";

dffeas A_ctrl_ld(
	.clk(clk_clk),
	.d(\M_ctrl_ld~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_ctrl_ld~q ),
	.prn(vcc));
defparam A_ctrl_ld.is_wysiwyg = "true";
defparam A_ctrl_ld.power_up = "low";

dffeas \A_slow_inst_result[0] (
	.clk(clk_clk),
	.d(\A_slow_inst_result_nxt[0]~0_combout ),
	.asdata(d_readdata[0]),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_ctrl_ld32~q ),
	.ena(\A_ctrl_ld~q ),
	.q(\A_slow_inst_result[0]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[0] .is_wysiwyg = "true";
defparam \A_slow_inst_result[0] .power_up = "low";

cyclonev_lcell_comb \D_ctrl_shift_right_arith~1 (
	.dataa(!\D_iw[14]~q ),
	.datab(!\D_ctrl_shift_right_arith~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_shift_right_arith~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_shift_right_arith~1 .extended_lut = "off";
defparam \D_ctrl_shift_right_arith~1 .lut_mask = 64'h7777777777777777;
defparam \D_ctrl_shift_right_arith~1 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_shift_right_arith~2 (
	.dataa(!\D_iw[15]~q ),
	.datab(!\D_iw[16]~q ),
	.datac(!\D_ctrl_shift_right_arith~1_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_shift_right_arith~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_shift_right_arith~2 .extended_lut = "off";
defparam \D_ctrl_shift_right_arith~2 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \D_ctrl_shift_right_arith~2 .shared_arith = "off";

dffeas E_ctrl_shift_right_arith(
	.clk(clk_clk),
	.d(\D_ctrl_shift_right_arith~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_ctrl_shift_right_arith~q ),
	.prn(vcc));
defparam E_ctrl_shift_right_arith.is_wysiwyg = "true";
defparam E_ctrl_shift_right_arith.power_up = "low";

cyclonev_lcell_comb \E_rot_fill_bit~0 (
	.dataa(!\E_src1[31]~q ),
	.datab(!\E_ctrl_shift_right_arith~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_fill_bit~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_fill_bit~0 .extended_lut = "off";
defparam \E_rot_fill_bit~0 .lut_mask = 64'h7777777777777777;
defparam \E_rot_fill_bit~0 .shared_arith = "off";

dffeas M_rot_fill_bit(
	.clk(clk_clk),
	.d(\E_rot_fill_bit~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_rot_fill_bit~q ),
	.prn(vcc));
defparam M_rot_fill_bit.is_wysiwyg = "true";
defparam M_rot_fill_bit.power_up = "low";

dffeas \M_alu_result[3] (
	.clk(clk_clk),
	.d(\E_alu_result[3]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_alu_result[3]~q ),
	.prn(vcc));
defparam \M_alu_result[3] .is_wysiwyg = "true";
defparam \M_alu_result[3] .power_up = "low";

dffeas \d_readdata_d1[3] (
	.clk(clk_clk),
	.d(d_readdata[3]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[3]~q ),
	.prn(vcc));
defparam \d_readdata_d1[3] .is_wysiwyg = "true";
defparam \d_readdata_d1[3] .power_up = "low";

dffeas \d_readdata_d1[19] (
	.clk(clk_clk),
	.d(d_readdata[19]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[19]~q ),
	.prn(vcc));
defparam \d_readdata_d1[19] .is_wysiwyg = "true";
defparam \d_readdata_d1[19] .power_up = "low";

dffeas \d_readdata_d1[11] (
	.clk(clk_clk),
	.d(d_readdata[11]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[11]~q ),
	.prn(vcc));
defparam \d_readdata_d1[11] .is_wysiwyg = "true";
defparam \d_readdata_d1[11] .power_up = "low";

dffeas \d_readdata_d1[27] (
	.clk(clk_clk),
	.d(d_readdata[27]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[27]~q ),
	.prn(vcc));
defparam \d_readdata_d1[27] .is_wysiwyg = "true";
defparam \d_readdata_d1[27] .power_up = "low";

cyclonev_lcell_comb \A_slow_inst_result_nxt[3]~3 (
	.dataa(!\d_readdata_d1[3]~q ),
	.datab(!\d_readdata_d1[19]~q ),
	.datac(!\d_readdata_d1[11]~q ),
	.datad(!\d_readdata_d1[27]~q ),
	.datae(!\A_ld_align_sh16~q ),
	.dataf(!\A_ld_align_sh8~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[3]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[3]~3 .extended_lut = "off";
defparam \A_slow_inst_result_nxt[3]~3 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_slow_inst_result_nxt[3]~3 .shared_arith = "off";

dffeas \A_slow_inst_result[3] (
	.clk(clk_clk),
	.d(\A_slow_inst_result_nxt[3]~3_combout ),
	.asdata(d_readdata[3]),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_ctrl_ld32~q ),
	.ena(\A_ctrl_ld~q ),
	.q(\A_slow_inst_result[3]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[3] .is_wysiwyg = "true";
defparam \A_slow_inst_result[3] .power_up = "low";

dffeas \M_alu_result[4] (
	.clk(clk_clk),
	.d(\E_alu_result[4]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_alu_result[4]~q ),
	.prn(vcc));
defparam \M_alu_result[4] .is_wysiwyg = "true";
defparam \M_alu_result[4] .power_up = "low";

dffeas \d_readdata_d1[4] (
	.clk(clk_clk),
	.d(d_readdata[4]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[4]~q ),
	.prn(vcc));
defparam \d_readdata_d1[4] .is_wysiwyg = "true";
defparam \d_readdata_d1[4] .power_up = "low";

dffeas \d_readdata_d1[20] (
	.clk(clk_clk),
	.d(d_readdata[20]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[20]~q ),
	.prn(vcc));
defparam \d_readdata_d1[20] .is_wysiwyg = "true";
defparam \d_readdata_d1[20] .power_up = "low";

dffeas \d_readdata_d1[12] (
	.clk(clk_clk),
	.d(d_readdata[12]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[12]~q ),
	.prn(vcc));
defparam \d_readdata_d1[12] .is_wysiwyg = "true";
defparam \d_readdata_d1[12] .power_up = "low";

dffeas \d_readdata_d1[28] (
	.clk(clk_clk),
	.d(d_readdata[28]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[28]~q ),
	.prn(vcc));
defparam \d_readdata_d1[28] .is_wysiwyg = "true";
defparam \d_readdata_d1[28] .power_up = "low";

cyclonev_lcell_comb \A_slow_inst_result_nxt[4]~4 (
	.dataa(!\d_readdata_d1[4]~q ),
	.datab(!\d_readdata_d1[20]~q ),
	.datac(!\d_readdata_d1[12]~q ),
	.datad(!\d_readdata_d1[28]~q ),
	.datae(!\A_ld_align_sh16~q ),
	.dataf(!\A_ld_align_sh8~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[4]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[4]~4 .extended_lut = "off";
defparam \A_slow_inst_result_nxt[4]~4 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_slow_inst_result_nxt[4]~4 .shared_arith = "off";

dffeas \A_slow_inst_result[4] (
	.clk(clk_clk),
	.d(\A_slow_inst_result_nxt[4]~4_combout ),
	.asdata(d_readdata[4]),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_ctrl_ld32~q ),
	.ena(\A_ctrl_ld~q ),
	.q(\A_slow_inst_result[4]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[4] .is_wysiwyg = "true";
defparam \A_slow_inst_result[4] .power_up = "low";

dffeas \M_alu_result[2] (
	.clk(clk_clk),
	.d(\E_alu_result[2]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_alu_result[2]~q ),
	.prn(vcc));
defparam \M_alu_result[2] .is_wysiwyg = "true";
defparam \M_alu_result[2] .power_up = "low";

dffeas \d_readdata_d1[2] (
	.clk(clk_clk),
	.d(d_readdata[2]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[2]~q ),
	.prn(vcc));
defparam \d_readdata_d1[2] .is_wysiwyg = "true";
defparam \d_readdata_d1[2] .power_up = "low";

dffeas \d_readdata_d1[18] (
	.clk(clk_clk),
	.d(d_readdata[18]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[18]~q ),
	.prn(vcc));
defparam \d_readdata_d1[18] .is_wysiwyg = "true";
defparam \d_readdata_d1[18] .power_up = "low";

dffeas \d_readdata_d1[10] (
	.clk(clk_clk),
	.d(d_readdata[10]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[10]~q ),
	.prn(vcc));
defparam \d_readdata_d1[10] .is_wysiwyg = "true";
defparam \d_readdata_d1[10] .power_up = "low";

dffeas \d_readdata_d1[26] (
	.clk(clk_clk),
	.d(d_readdata[26]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[26]~q ),
	.prn(vcc));
defparam \d_readdata_d1[26] .is_wysiwyg = "true";
defparam \d_readdata_d1[26] .power_up = "low";

cyclonev_lcell_comb \A_slow_inst_result_nxt[2]~2 (
	.dataa(!\d_readdata_d1[2]~q ),
	.datab(!\d_readdata_d1[18]~q ),
	.datac(!\d_readdata_d1[10]~q ),
	.datad(!\d_readdata_d1[26]~q ),
	.datae(!\A_ld_align_sh16~q ),
	.dataf(!\A_ld_align_sh8~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[2]~2 .extended_lut = "off";
defparam \A_slow_inst_result_nxt[2]~2 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_slow_inst_result_nxt[2]~2 .shared_arith = "off";

dffeas \A_slow_inst_result[2] (
	.clk(clk_clk),
	.d(\A_slow_inst_result_nxt[2]~2_combout ),
	.asdata(d_readdata[2]),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_ctrl_ld32~q ),
	.ena(\A_ctrl_ld~q ),
	.q(\A_slow_inst_result[2]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[2] .is_wysiwyg = "true";
defparam \A_slow_inst_result[2] .power_up = "low";

dffeas E_ctrl_shift_rot_right(
	.clk(clk_clk),
	.d(\D_ctrl_shift_right_arith~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_ctrl_shift_rot_right~q ),
	.prn(vcc));
defparam E_ctrl_shift_rot_right.is_wysiwyg = "true";
defparam E_ctrl_shift_rot_right.power_up = "low";

cyclonev_lcell_comb \E_rot_mask[2]~2 (
	.dataa(!\E_src2[2]~q ),
	.datab(!\E_src2[1]~q ),
	.datac(!\E_src2[0]~q ),
	.datad(!\E_ctrl_shift_rot_right~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_mask[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_mask[2]~2 .extended_lut = "off";
defparam \E_rot_mask[2]~2 .lut_mask = 64'hFF7FFF7FFF7FFF7F;
defparam \E_rot_mask[2]~2 .shared_arith = "off";

dffeas \M_rot_mask[2] (
	.clk(clk_clk),
	.d(\E_rot_mask[2]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_rot_mask[2]~q ),
	.prn(vcc));
defparam \M_rot_mask[2] .is_wysiwyg = "true";
defparam \M_rot_mask[2] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[0]~7 (
	.dataa(!\D_ctrl_b_is_dst~q ),
	.datab(!\A_regnum_b_cmp_D~q ),
	.datac(!\M_regnum_b_cmp_D~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[0]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[0]~7 .extended_lut = "off";
defparam \D_src2_reg[0]~7 .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \D_src2_reg[0]~7 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[0]~8 (
	.dataa(!\D_ctrl_b_is_dst~q ),
	.datab(!\W_regnum_b_cmp_D~q ),
	.datac(!\A_regnum_b_cmp_D~q ),
	.datad(!\M_regnum_b_cmp_D~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[0]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[0]~8 .extended_lut = "off";
defparam \D_src2_reg[0]~8 .lut_mask = 64'hFFBFFFBFFFBFFFBF;
defparam \D_src2_reg[0]~8 .shared_arith = "off";

dffeas M_ctrl_ld8_ld16(
	.clk(clk_clk),
	.d(\Equal212~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_ctrl_ld8_ld16~q ),
	.prn(vcc));
defparam M_ctrl_ld8_ld16.is_wysiwyg = "true";
defparam M_ctrl_ld8_ld16.power_up = "low";

cyclonev_lcell_comb M_ld_align_byte2_byte3_fill(
	.dataa(!\M_exc_any~combout ),
	.datab(!\M_ctrl_ld8_ld16~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_ld_align_byte2_byte3_fill~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam M_ld_align_byte2_byte3_fill.extended_lut = "off";
defparam M_ld_align_byte2_byte3_fill.lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam M_ld_align_byte2_byte3_fill.shared_arith = "off";

dffeas A_ld_align_byte2_byte3_fill(
	.clk(clk_clk),
	.d(\M_ld_align_byte2_byte3_fill~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_ld_align_byte2_byte3_fill~q ),
	.prn(vcc));
defparam A_ld_align_byte2_byte3_fill.is_wysiwyg = "true";
defparam A_ld_align_byte2_byte3_fill.power_up = "low";

dffeas \d_readdata_d1[22] (
	.clk(clk_clk),
	.d(d_readdata[22]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[22]~q ),
	.prn(vcc));
defparam \d_readdata_d1[22] .is_wysiwyg = "true";
defparam \d_readdata_d1[22] .power_up = "low";

cyclonev_lcell_comb \A_slow_inst_result_nxt[22]~35 (
	.dataa(!\A_ctrl_ld32~q ),
	.datab(!\d_readdata_d1[22]~q ),
	.datac(!read_latency_shift_reg_01),
	.datad(!src0_valid),
	.datae(!av_readdata_pre_22),
	.dataf(!av_readdata_pre_221),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[22]~35_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[22]~35 .extended_lut = "off";
defparam \A_slow_inst_result_nxt[22]~35 .lut_mask = 64'h27FFFFFFFFFFFFFF;
defparam \A_slow_inst_result_nxt[22]~35 .shared_arith = "off";

cyclonev_lcell_comb \A_slow_inst_result_nxt[22]~8 (
	.dataa(!\A_ctrl_ld32~q ),
	.datab(!\A_ld_align_byte2_byte3_fill~q ),
	.datac(!\A_slow_ld_data_fill_bit~0_combout ),
	.datad(!src0_valid1),
	.datae(!q_a_22),
	.dataf(!\A_slow_inst_result_nxt[22]~35_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[22]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[22]~8 .extended_lut = "off";
defparam \A_slow_inst_result_nxt[22]~8 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \A_slow_inst_result_nxt[22]~8 .shared_arith = "off";

dffeas \A_slow_inst_result[22] (
	.clk(clk_clk),
	.d(\A_slow_inst_result_nxt[22]~8_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_ctrl_ld~q ),
	.q(\A_slow_inst_result[22]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[22] .is_wysiwyg = "true";
defparam \A_slow_inst_result[22] .power_up = "low";

cyclonev_lcell_comb \E_rot_mask[6]~6 (
	.dataa(!\E_src2[2]~q ),
	.datab(!\E_src2[1]~q ),
	.datac(!\E_src2[0]~q ),
	.datad(!\E_ctrl_shift_rot_right~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_mask[6]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_mask[6]~6 .extended_lut = "off";
defparam \E_rot_mask[6]~6 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \E_rot_mask[6]~6 .shared_arith = "off";

dffeas \M_rot_mask[6] (
	.clk(clk_clk),
	.d(\E_rot_mask[6]~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_rot_mask[6]~q ),
	.prn(vcc));
defparam \M_rot_mask[6] .is_wysiwyg = "true";
defparam \M_rot_mask[6] .power_up = "low";

cyclonev_lcell_comb \D_ctrl_rot~0 (
	.dataa(!\D_iw[15]~q ),
	.datab(!\D_ctrl_shift_right_arith~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_rot~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_rot~0 .extended_lut = "off";
defparam \D_ctrl_rot~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \D_ctrl_rot~0 .shared_arith = "off";

dffeas E_ctrl_rot(
	.clk(clk_clk),
	.d(\D_ctrl_rot~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_ctrl_rot~q ),
	.prn(vcc));
defparam E_ctrl_rot.is_wysiwyg = "true";
defparam E_ctrl_rot.power_up = "low";

cyclonev_lcell_comb \D_ctrl_shift_rot_left~0 (
	.dataa(!\D_iw[14]~q ),
	.datab(!\D_ctrl_shift_right_arith~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_shift_rot_left~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_shift_rot_left~0 .extended_lut = "off";
defparam \D_ctrl_shift_rot_left~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \D_ctrl_shift_rot_left~0 .shared_arith = "off";

dffeas E_ctrl_shift_rot_left(
	.clk(clk_clk),
	.d(\D_ctrl_shift_rot_left~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_ctrl_shift_rot_left~q ),
	.prn(vcc));
defparam E_ctrl_shift_rot_left.is_wysiwyg = "true";
defparam E_ctrl_shift_rot_left.power_up = "low";

cyclonev_lcell_comb \E_rot_pass2~0 (
	.dataa(!\E_src2[3]~q ),
	.datab(!\E_src2[4]~q ),
	.datac(!\E_ctrl_rot~q ),
	.datad(!\E_ctrl_shift_rot_right~q ),
	.datae(!\E_ctrl_shift_rot_left~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_pass2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_pass2~0 .extended_lut = "off";
defparam \E_rot_pass2~0 .lut_mask = 64'hEFFFFFFFEFFFFFFF;
defparam \E_rot_pass2~0 .shared_arith = "off";

dffeas M_rot_pass2(
	.clk(clk_clk),
	.d(\E_rot_pass2~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_rot_pass2~q ),
	.prn(vcc));
defparam M_rot_pass2.is_wysiwyg = "true";
defparam M_rot_pass2.power_up = "low";

cyclonev_lcell_comb \E_rot_sel_fill2~0 (
	.dataa(!\E_src2[3]~q ),
	.datab(!\E_src2[4]~q ),
	.datac(!\E_ctrl_shift_rot_right~q ),
	.datad(!\E_ctrl_shift_rot_left~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_sel_fill2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_sel_fill2~0 .extended_lut = "off";
defparam \E_rot_sel_fill2~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \E_rot_sel_fill2~0 .shared_arith = "off";

dffeas M_rot_sel_fill2(
	.clk(clk_clk),
	.d(\E_rot_sel_fill2~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_rot_sel_fill2~q ),
	.prn(vcc));
defparam M_rot_sel_fill2.is_wysiwyg = "true";
defparam M_rot_sel_fill2.power_up = "low";

cyclonev_lcell_comb \A_slow_inst_result_nxt[18]~32 (
	.dataa(!\A_ctrl_ld32~q ),
	.datab(!\A_ld_align_byte2_byte3_fill~q ),
	.datac(!src0_valid),
	.datad(!av_readdata_pre_18),
	.datae(!src_payload10),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[18]~32_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[18]~32 .extended_lut = "off";
defparam \A_slow_inst_result_nxt[18]~32 .lut_mask = 64'hFFD8FFFFFFD8FFFF;
defparam \A_slow_inst_result_nxt[18]~32 .shared_arith = "off";

cyclonev_lcell_comb \A_slow_inst_result_nxt[18]~21 (
	.dataa(!\A_ctrl_ld32~q ),
	.datab(!\d_readdata_d1[18]~q ),
	.datac(!\A_slow_ld_data_fill_bit~0_combout ),
	.datad(!src0_valid1),
	.datae(!q_a_18),
	.dataf(!\A_slow_inst_result_nxt[18]~32_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[18]~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[18]~21 .extended_lut = "off";
defparam \A_slow_inst_result_nxt[18]~21 .lut_mask = 64'h7FFFFFFFBFFFFFFF;
defparam \A_slow_inst_result_nxt[18]~21 .shared_arith = "off";

dffeas \A_slow_inst_result[18] (
	.clk(clk_clk),
	.d(\A_slow_inst_result_nxt[18]~21_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_ctrl_ld~q ),
	.q(\A_slow_inst_result[18]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[18] .is_wysiwyg = "true";
defparam \A_slow_inst_result[18] .power_up = "low";

cyclonev_lcell_comb \M_ld_align_byte1_fill~0 (
	.dataa(!\M_exc_any~combout ),
	.datab(!\M_ctrl_ld8~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_ld_align_byte1_fill~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_ld_align_byte1_fill~0 .extended_lut = "off";
defparam \M_ld_align_byte1_fill~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \M_ld_align_byte1_fill~0 .shared_arith = "off";

dffeas A_ld_align_byte1_fill(
	.clk(clk_clk),
	.d(\M_ld_align_byte1_fill~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_ld_align_byte1_fill~q ),
	.prn(vcc));
defparam A_ld_align_byte1_fill.is_wysiwyg = "true";
defparam A_ld_align_byte1_fill.power_up = "low";

cyclonev_lcell_comb \A_slow_inst_result[9]~1 (
	.dataa(!\A_ctrl_ld32~q ),
	.datab(!\A_ld_align_byte1_fill~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result[9]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result[9]~1 .extended_lut = "off";
defparam \A_slow_inst_result[9]~1 .lut_mask = 64'h7777777777777777;
defparam \A_slow_inst_result[9]~1 .shared_arith = "off";

dffeas \d_readdata_d1[14] (
	.clk(clk_clk),
	.d(d_readdata[14]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[14]~q ),
	.prn(vcc));
defparam \d_readdata_d1[14] .is_wysiwyg = "true";
defparam \d_readdata_d1[14] .power_up = "low";

dffeas \d_readdata_d1[30] (
	.clk(clk_clk),
	.d(d_readdata[30]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[30]~q ),
	.prn(vcc));
defparam \d_readdata_d1[30] .is_wysiwyg = "true";
defparam \d_readdata_d1[30] .power_up = "low";

cyclonev_lcell_comb \A_slow_inst_result[9]~0 (
	.dataa(!\A_ctrl_ld32~q ),
	.datab(!\A_ld_align_sh16~q ),
	.datac(!\A_ld_align_byte1_fill~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result[9]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result[9]~0 .extended_lut = "off";
defparam \A_slow_inst_result[9]~0 .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \A_slow_inst_result[9]~0 .shared_arith = "off";

cyclonev_lcell_comb \A_slow_inst_result_nxt[14]~46 (
	.dataa(!\d_readdata_d1[14]~q ),
	.datab(!\d_readdata_d1[30]~q ),
	.datac(!\A_slow_inst_result[9]~0_combout ),
	.datad(!\A_slow_inst_result[9]~1_combout ),
	.datae(!src0_valid),
	.dataf(!av_readdata_pre_14),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[14]~46_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[14]~46 .extended_lut = "off";
defparam \A_slow_inst_result_nxt[14]~46 .lut_mask = 64'h7FF7FFFFFFFFFFFF;
defparam \A_slow_inst_result_nxt[14]~46 .shared_arith = "off";

cyclonev_lcell_comb \A_slow_inst_result_nxt[14]~48 (
	.dataa(!\A_slow_inst_result[9]~1_combout ),
	.datab(!\A_slow_inst_result_nxt[14]~46_combout ),
	.datac(!\A_slow_ld_data_fill_bit~0_combout ),
	.datad(!src_payload15),
	.datae(!\A_slow_inst_result[9]~0_combout ),
	.dataf(!q_a_14),
	.datag(!src0_valid1),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[14]~48_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[14]~48 .extended_lut = "on";
defparam \A_slow_inst_result_nxt[14]~48 .lut_mask = 64'hFFD8FFD8FFD8FFD8;
defparam \A_slow_inst_result_nxt[14]~48 .shared_arith = "off";

dffeas \A_slow_inst_result[14] (
	.clk(clk_clk),
	.d(\A_slow_inst_result_nxt[14]~48_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_ctrl_ld~q ),
	.q(\A_slow_inst_result[14]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[14] .is_wysiwyg = "true";
defparam \A_slow_inst_result[14] .power_up = "low";

cyclonev_lcell_comb \E_rot_pass1~0 (
	.dataa(!\E_src2[3]~q ),
	.datab(!\E_src2[4]~q ),
	.datac(!\E_ctrl_rot~q ),
	.datad(!\E_ctrl_shift_rot_right~q ),
	.datae(!\E_ctrl_shift_rot_left~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_pass1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_pass1~0 .extended_lut = "off";
defparam \E_rot_pass1~0 .lut_mask = 64'hEFFFFFFFEFFFFFFF;
defparam \E_rot_pass1~0 .shared_arith = "off";

dffeas M_rot_pass1(
	.clk(clk_clk),
	.d(\E_rot_pass1~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_rot_pass1~q ),
	.prn(vcc));
defparam M_rot_pass1.is_wysiwyg = "true";
defparam M_rot_pass1.power_up = "low";

cyclonev_lcell_comb \E_rot_sel_fill1~0 (
	.dataa(!\E_src2[3]~q ),
	.datab(!\E_src2[4]~q ),
	.datac(!\E_ctrl_shift_rot_right~q ),
	.datad(!\E_ctrl_shift_rot_left~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_sel_fill1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_sel_fill1~0 .extended_lut = "off";
defparam \E_rot_sel_fill1~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \E_rot_sel_fill1~0 .shared_arith = "off";

dffeas M_rot_sel_fill1(
	.clk(clk_clk),
	.d(\E_rot_sel_fill1~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_rot_sel_fill1~q ),
	.prn(vcc));
defparam M_rot_sel_fill1.is_wysiwyg = "true";
defparam M_rot_sel_fill1.power_up = "low";

cyclonev_lcell_comb \A_slow_inst_result_nxt[10]~42 (
	.dataa(!\d_readdata_d1[10]~q ),
	.datab(!\d_readdata_d1[26]~q ),
	.datac(!\A_slow_inst_result[9]~0_combout ),
	.datad(!\A_slow_inst_result[9]~1_combout ),
	.datae(!src0_valid),
	.dataf(!av_readdata_pre_10),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[10]~42_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[10]~42 .extended_lut = "off";
defparam \A_slow_inst_result_nxt[10]~42 .lut_mask = 64'h7FF7FFFFFFFFFFFF;
defparam \A_slow_inst_result_nxt[10]~42 .shared_arith = "off";

cyclonev_lcell_comb \A_slow_inst_result_nxt[10]~72 (
	.dataa(!\A_slow_inst_result_nxt[10]~42_combout ),
	.datab(!q_a_10),
	.datac(!\A_slow_ld_data_fill_bit~0_combout ),
	.datad(!src0_valid1),
	.datae(!\A_slow_inst_result[9]~0_combout ),
	.dataf(!\A_slow_inst_result[9]~1_combout ),
	.datag(!src_payload6),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[10]~72_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[10]~72 .extended_lut = "on";
defparam \A_slow_inst_result_nxt[10]~72 .lut_mask = 64'hFFD8FFD8FFD8FFD8;
defparam \A_slow_inst_result_nxt[10]~72 .shared_arith = "off";

dffeas \A_slow_inst_result[10] (
	.clk(clk_clk),
	.d(\A_slow_inst_result_nxt[10]~72_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_ctrl_ld~q ),
	.q(\A_slow_inst_result[10]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[10] .is_wysiwyg = "true";
defparam \A_slow_inst_result[10] .power_up = "low";

dffeas \d_readdata_d1[6] (
	.clk(clk_clk),
	.d(d_readdata[6]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[6]~q ),
	.prn(vcc));
defparam \d_readdata_d1[6] .is_wysiwyg = "true";
defparam \d_readdata_d1[6] .power_up = "low";

cyclonev_lcell_comb \A_slow_inst_result_nxt[6]~6 (
	.dataa(!\d_readdata_d1[6]~q ),
	.datab(!\d_readdata_d1[22]~q ),
	.datac(!\d_readdata_d1[14]~q ),
	.datad(!\d_readdata_d1[30]~q ),
	.datae(!\A_ld_align_sh16~q ),
	.dataf(!\A_ld_align_sh8~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[6]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[6]~6 .extended_lut = "off";
defparam \A_slow_inst_result_nxt[6]~6 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_slow_inst_result_nxt[6]~6 .shared_arith = "off";

dffeas \A_slow_inst_result[6] (
	.clk(clk_clk),
	.d(\A_slow_inst_result_nxt[6]~6_combout ),
	.asdata(d_readdata[6]),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_ctrl_ld32~q ),
	.ena(\A_ctrl_ld~q ),
	.q(\A_slow_inst_result[6]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[6] .is_wysiwyg = "true";
defparam \A_slow_inst_result[6] .power_up = "low";

dffeas \E_compare_op[0] (
	.clk(clk_clk),
	.d(\D_logic_op_raw[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_compare_op[0]~q ),
	.prn(vcc));
defparam \E_compare_op[0] .is_wysiwyg = "true";
defparam \E_compare_op[0] .power_up = "low";

cyclonev_lcell_comb \E_logic_result[3]~0 (
	.dataa(!\E_src2[3]~q ),
	.datab(!\E_src1[3]~q ),
	.datac(!\E_logic_op[1]~q ),
	.datad(!\E_logic_op[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[3]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[3]~0 .extended_lut = "off";
defparam \E_logic_result[3]~0 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[3]~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal316~0 (
	.dataa(!\E_src2[0]~q ),
	.datab(!\E_src1[0]~q ),
	.datac(!\E_src2[25]~q ),
	.datad(!\E_src1[25]~q ),
	.datae(!\E_logic_op[1]~q ),
	.dataf(!\E_logic_op[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal316~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal316~0 .extended_lut = "off";
defparam \Equal316~0 .lut_mask = 64'h6996966996696996;
defparam \Equal316~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal316~1 (
	.dataa(!\E_src2[2]~q ),
	.datab(!\E_src1[2]~q ),
	.datac(!\E_src2[31]~q ),
	.datad(!\E_src1[31]~q ),
	.datae(!\E_logic_op[1]~q ),
	.dataf(!\E_logic_op[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal316~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal316~1 .extended_lut = "off";
defparam \Equal316~1 .lut_mask = 64'h6996966996696996;
defparam \Equal316~1 .shared_arith = "off";

cyclonev_lcell_comb \Equal316~2 (
	.dataa(!\E_logic_result[3]~0_combout ),
	.datab(!\E_logic_result[22]~1_combout ),
	.datac(!\E_logic_result[23]~2_combout ),
	.datad(!\E_logic_result[24]~3_combout ),
	.datae(!\Equal316~0_combout ),
	.dataf(!\Equal316~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal316~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal316~2 .extended_lut = "off";
defparam \Equal316~2 .lut_mask = 64'hFFFEFFFFFFFFFFFF;
defparam \Equal316~2 .shared_arith = "off";

dffeas \d_readdata_d1[7] (
	.clk(clk_clk),
	.d(d_readdata[7]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[7]~q ),
	.prn(vcc));
defparam \d_readdata_d1[7] .is_wysiwyg = "true";
defparam \d_readdata_d1[7] .power_up = "low";

dffeas \d_readdata_d1[23] (
	.clk(clk_clk),
	.d(d_readdata[23]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[23]~q ),
	.prn(vcc));
defparam \d_readdata_d1[23] .is_wysiwyg = "true";
defparam \d_readdata_d1[23] .power_up = "low";

dffeas \d_readdata_d1[15] (
	.clk(clk_clk),
	.d(d_readdata[15]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[15]~q ),
	.prn(vcc));
defparam \d_readdata_d1[15] .is_wysiwyg = "true";
defparam \d_readdata_d1[15] .power_up = "low";

cyclonev_lcell_comb \A_slow_inst_result_nxt[7]~7 (
	.dataa(!\d_readdata_d1[7]~q ),
	.datab(!\d_readdata_d1[23]~q ),
	.datac(!\d_readdata_d1[15]~q ),
	.datad(!\d_readdata_d1[31]~q ),
	.datae(!\A_ld_align_sh16~q ),
	.dataf(!\A_ld_align_sh8~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[7]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[7]~7 .extended_lut = "off";
defparam \A_slow_inst_result_nxt[7]~7 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_slow_inst_result_nxt[7]~7 .shared_arith = "off";

dffeas \A_slow_inst_result[7] (
	.clk(clk_clk),
	.d(\A_slow_inst_result_nxt[7]~7_combout ),
	.asdata(d_readdata[7]),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_ctrl_ld32~q ),
	.ena(\A_ctrl_ld~q ),
	.q(\A_slow_inst_result[7]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[7] .is_wysiwyg = "true";
defparam \A_slow_inst_result[7] .power_up = "low";

cyclonev_lcell_comb \E_rot_mask[7]~7 (
	.dataa(!\E_src2[2]~q ),
	.datab(!\E_src2[1]~q ),
	.datac(!\E_src2[0]~q ),
	.datad(!\E_ctrl_shift_rot_right~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_mask[7]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_mask[7]~7 .extended_lut = "off";
defparam \E_rot_mask[7]~7 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \E_rot_mask[7]~7 .shared_arith = "off";

dffeas \M_rot_mask[7] (
	.clk(clk_clk),
	.d(\E_rot_mask[7]~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_rot_mask[7]~q ),
	.prn(vcc));
defparam \M_rot_mask[7] .is_wysiwyg = "true";
defparam \M_rot_mask[7] .power_up = "low";

cyclonev_lcell_comb \Add10~0 (
	.dataa(!\E_src2[1]~q ),
	.datab(!\E_src2[0]~q ),
	.datac(!\E_ctrl_shift_rot_right~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add10~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add10~0 .extended_lut = "off";
defparam \Add10~0 .lut_mask = 64'h9696969696969696;
defparam \Add10~0 .shared_arith = "off";

cyclonev_lcell_comb \E_rot_step1[3]~25 (
	.dataa(!\E_src1[3]~q ),
	.datab(!\E_src1[2]~q ),
	.datac(!\E_src1[1]~q ),
	.datad(!\E_src1[0]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add10~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[3]~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[3]~25 .extended_lut = "off";
defparam \E_rot_step1[3]~25 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[3]~25 .shared_arith = "off";

dffeas \d_readdata_d1[5] (
	.clk(clk_clk),
	.d(d_readdata[5]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[5]~q ),
	.prn(vcc));
defparam \d_readdata_d1[5] .is_wysiwyg = "true";
defparam \d_readdata_d1[5] .power_up = "low";

dffeas \d_readdata_d1[21] (
	.clk(clk_clk),
	.d(d_readdata[21]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[21]~q ),
	.prn(vcc));
defparam \d_readdata_d1[21] .is_wysiwyg = "true";
defparam \d_readdata_d1[21] .power_up = "low";

dffeas \d_readdata_d1[13] (
	.clk(clk_clk),
	.d(d_readdata[13]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[13]~q ),
	.prn(vcc));
defparam \d_readdata_d1[13] .is_wysiwyg = "true";
defparam \d_readdata_d1[13] .power_up = "low";

dffeas \d_readdata_d1[29] (
	.clk(clk_clk),
	.d(d_readdata[29]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[29]~q ),
	.prn(vcc));
defparam \d_readdata_d1[29] .is_wysiwyg = "true";
defparam \d_readdata_d1[29] .power_up = "low";

cyclonev_lcell_comb \A_slow_inst_result_nxt[5]~5 (
	.dataa(!\d_readdata_d1[5]~q ),
	.datab(!\d_readdata_d1[21]~q ),
	.datac(!\d_readdata_d1[13]~q ),
	.datad(!\d_readdata_d1[29]~q ),
	.datae(!\A_ld_align_sh16~q ),
	.dataf(!\A_ld_align_sh8~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[5]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[5]~5 .extended_lut = "off";
defparam \A_slow_inst_result_nxt[5]~5 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_slow_inst_result_nxt[5]~5 .shared_arith = "off";

dffeas \A_slow_inst_result[5] (
	.clk(clk_clk),
	.d(\A_slow_inst_result_nxt[5]~5_combout ),
	.asdata(d_readdata[5]),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_ctrl_ld32~q ),
	.ena(\A_ctrl_ld~q ),
	.q(\A_slow_inst_result[5]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[5] .is_wysiwyg = "true";
defparam \A_slow_inst_result[5] .power_up = "low";

cyclonev_lcell_comb \E_rot_mask[5]~5 (
	.dataa(!\E_src2[2]~q ),
	.datab(!\E_src2[1]~q ),
	.datac(!\E_src2[0]~q ),
	.datad(!\E_ctrl_shift_rot_right~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_mask[5]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_mask[5]~5 .extended_lut = "off";
defparam \E_rot_mask[5]~5 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \E_rot_mask[5]~5 .shared_arith = "off";

dffeas \M_rot_mask[5] (
	.clk(clk_clk),
	.d(\E_rot_mask[5]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_rot_mask[5]~q ),
	.prn(vcc));
defparam \M_rot_mask[5] .is_wysiwyg = "true";
defparam \M_rot_mask[5] .power_up = "low";

cyclonev_lcell_comb \E_rot_step1[1]~9 (
	.dataa(!\E_src1[1]~q ),
	.datab(!\E_src1[0]~q ),
	.datac(!\E_src1[31]~q ),
	.datad(!\E_src1[30]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add10~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[1]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[1]~9 .extended_lut = "off";
defparam \E_rot_step1[1]~9 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[1]~9 .shared_arith = "off";

cyclonev_lcell_comb \Add9~134 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\Add9~134_cout ),
	.shareout());
defparam \Add9~134 .extended_lut = "off";
defparam \Add9~134 .lut_mask = 64'h0000000000005555;
defparam \Add9~134 .shared_arith = "off";

cyclonev_lcell_comb \Add9~65 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[0]~q ),
	.datae(gnd),
	.dataf(!\E_src1[0]~q ),
	.datag(gnd),
	.cin(\Add9~134_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~65_sumout ),
	.cout(\Add9~66 ),
	.shareout());
defparam \Add9~65 .extended_lut = "off";
defparam \Add9~65 .lut_mask = 64'h0000FF00000055AA;
defparam \Add9~65 .shared_arith = "off";

cyclonev_lcell_comb \Add9~69 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[1]~q ),
	.datae(gnd),
	.dataf(!\E_src1[1]~q ),
	.datag(gnd),
	.cin(\Add9~66 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~69_sumout ),
	.cout(\Add9~70 ),
	.shareout());
defparam \Add9~69 .extended_lut = "off";
defparam \Add9~69 .lut_mask = 64'h0000FF00000055AA;
defparam \Add9~69 .shared_arith = "off";

cyclonev_lcell_comb \Add9~57 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[2]~q ),
	.datae(gnd),
	.dataf(!\E_src1[2]~q ),
	.datag(gnd),
	.cin(\Add9~70 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~57_sumout ),
	.cout(\Add9~58 ),
	.shareout());
defparam \Add9~57 .extended_lut = "off";
defparam \Add9~57 .lut_mask = 64'h0000FF00000055AA;
defparam \Add9~57 .shared_arith = "off";

cyclonev_lcell_comb \Add9~53 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[3]~q ),
	.datae(gnd),
	.dataf(!\E_src1[3]~q ),
	.datag(gnd),
	.cin(\Add9~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~53_sumout ),
	.cout(\Add9~54 ),
	.shareout());
defparam \Add9~53 .extended_lut = "off";
defparam \Add9~53 .lut_mask = 64'h0000FF00000055AA;
defparam \Add9~53 .shared_arith = "off";

cyclonev_lcell_comb \Add9~1 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[4]~q ),
	.datae(gnd),
	.dataf(!\E_src1[4]~q ),
	.datag(gnd),
	.cin(\Add9~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~1_sumout ),
	.cout(\Add9~2 ),
	.shareout());
defparam \Add9~1 .extended_lut = "off";
defparam \Add9~1 .lut_mask = 64'h0000FF00000055AA;
defparam \Add9~1 .shared_arith = "off";

cyclonev_lcell_comb \Add9~5 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[5]~q ),
	.datae(gnd),
	.dataf(!\E_src1[5]~q ),
	.datag(gnd),
	.cin(\Add9~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~5_sumout ),
	.cout(\Add9~6 ),
	.shareout());
defparam \Add9~5 .extended_lut = "off";
defparam \Add9~5 .lut_mask = 64'h0000FF00000055AA;
defparam \Add9~5 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result~4 (
	.dataa(!\E_src2[5]~q ),
	.datab(!\E_src1[5]~q ),
	.datac(!\E_logic_op[1]~q ),
	.datad(!\E_logic_op[0]~q ),
	.datae(!\E_ctrl_logic~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result~4 .extended_lut = "off";
defparam \E_alu_result~4 .lut_mask = 64'h6996FFFF6996FFFF;
defparam \E_alu_result~4 .shared_arith = "off";

dffeas \D_pc[3] (
	.clk(clk_clk),
	.d(\F_pc[3]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_pc[3]~q ),
	.prn(vcc));
defparam \D_pc[3] .is_wysiwyg = "true";
defparam \D_pc[3] .power_up = "low";

dffeas \D_iw[9] (
	.clk(clk_clk),
	.d(\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[9] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_iw[9]~q ),
	.prn(vcc));
defparam \D_iw[9] .is_wysiwyg = "true";
defparam \D_iw[9] .power_up = "low";

cyclonev_lcell_comb \Equal95~6 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[1]~q ),
	.datac(!\D_iw[2]~q ),
	.datad(!\D_iw[3]~q ),
	.datae(!\D_iw[4]~q ),
	.dataf(!\D_iw[5]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal95~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal95~6 .extended_lut = "off";
defparam \Equal95~6 .lut_mask = 64'hFFFFFFFFFFFFFFFD;
defparam \Equal95~6 .shared_arith = "off";

cyclonev_lcell_comb \F_ctrl_br~0 (
	.dataa(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[1] ),
	.datab(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[0] ),
	.datac(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[2] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ctrl_br~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ctrl_br~0 .extended_lut = "off";
defparam \F_ctrl_br~0 .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \F_ctrl_br~0 .shared_arith = "off";

dffeas D_ctrl_br(
	.clk(clk_clk),
	.d(\F_ctrl_br~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_ctrl_br~q ),
	.prn(vcc));
defparam D_ctrl_br.is_wysiwyg = "true";
defparam D_ctrl_br.power_up = "low";

dffeas \D_bht_data[1] (
	.clk(clk_clk),
	.d(\first_nios2_system_cpu_cpu_bht|the_altsyncram|auto_generated|q_b[1] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_bht_data[1]~q ),
	.prn(vcc));
defparam \D_bht_data[1] .is_wysiwyg = "true";
defparam \D_bht_data[1] .power_up = "low";

cyclonev_lcell_comb \F_ctrl_br_uncond~0 (
	.dataa(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[1] ),
	.datab(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[0] ),
	.datac(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[3] ),
	.datad(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[4] ),
	.datae(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[5] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ctrl_br_uncond~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ctrl_br_uncond~0 .extended_lut = "off";
defparam \F_ctrl_br_uncond~0 .lut_mask = 64'hFFFFFFFDFFFFFFFD;
defparam \F_ctrl_br_uncond~0 .shared_arith = "off";

dffeas D_ctrl_br_uncond(
	.clk(clk_clk),
	.d(\F_ctrl_br_uncond~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_ctrl_br_uncond~q ),
	.prn(vcc));
defparam D_ctrl_br_uncond.is_wysiwyg = "true";
defparam D_ctrl_br_uncond.power_up = "low";

cyclonev_lcell_comb \D_br_pred_taken~0 (
	.dataa(!\D_ctrl_br~q ),
	.datab(!\D_bht_data[1]~q ),
	.datac(!\D_ctrl_br_uncond~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_br_pred_taken~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_br_pred_taken~0 .extended_lut = "off";
defparam \D_br_pred_taken~0 .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \D_br_pred_taken~0 .shared_arith = "off";

cyclonev_lcell_comb \F_older_non_sequential~0 (
	.dataa(!\D_iw[16]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[11]~q ),
	.datad(!\Equal95~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_older_non_sequential~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_older_non_sequential~0 .extended_lut = "off";
defparam \F_older_non_sequential~0 .lut_mask = 64'hEFFFEFFFEFFFEFFF;
defparam \F_older_non_sequential~0 .shared_arith = "off";

cyclonev_lcell_comb \E_ctrl_jmp_indirect_nxt~0 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[16]~q ),
	.datad(!\Equal95~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_ctrl_jmp_indirect_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_ctrl_jmp_indirect_nxt~0 .extended_lut = "off";
defparam \E_ctrl_jmp_indirect_nxt~0 .lut_mask = 64'hFDFFFDFFFDFFFDFF;
defparam \E_ctrl_jmp_indirect_nxt~0 .shared_arith = "off";

cyclonev_lcell_comb \E_valid_jmp_indirect~0 (
	.dataa(!\E_ctrl_jmp_indirect_nxt~0_combout ),
	.datab(!\D_valid~combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_valid_jmp_indirect~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_valid_jmp_indirect~0 .extended_lut = "off";
defparam \E_valid_jmp_indirect~0 .lut_mask = 64'h7777777777777777;
defparam \E_valid_jmp_indirect~0 .shared_arith = "off";

dffeas E_valid_jmp_indirect(
	.clk(clk_clk),
	.d(\E_valid_jmp_indirect~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_valid_jmp_indirect~q ),
	.prn(vcc));
defparam E_valid_jmp_indirect.is_wysiwyg = "true";
defparam E_valid_jmp_indirect.power_up = "low";

dffeas \D_pc[2] (
	.clk(clk_clk),
	.d(\F_pc[2]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_pc[2]~q ),
	.prn(vcc));
defparam \D_pc[2] .is_wysiwyg = "true";
defparam \D_pc[2] .power_up = "low";

dffeas \D_pc[1] (
	.clk(clk_clk),
	.d(\F_pc[1]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_pc[1]~q ),
	.prn(vcc));
defparam \D_pc[1] .is_wysiwyg = "true";
defparam \D_pc[1] .power_up = "low";

dffeas \D_pc[0] (
	.clk(clk_clk),
	.d(\F_pc[0]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_pc[0]~q ),
	.prn(vcc));
defparam \D_pc[0] .is_wysiwyg = "true";
defparam \D_pc[0] .power_up = "low";

cyclonev_lcell_comb \Add3~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\F_pc[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~1_sumout ),
	.cout(\Add3~2 ),
	.shareout());
defparam \Add3~1 .extended_lut = "off";
defparam \Add3~1 .lut_mask = 64'h00000000000000FF;
defparam \Add3~1 .shared_arith = "off";

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[8] ),
	.datae(gnd),
	.dataf(!\Add3~1_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(\Add0~2 ),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~1 .shared_arith = "off";

dffeas \D_br_taken_waddr_partial[0] (
	.clk(clk_clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_br_taken_waddr_partial[0]~q ),
	.prn(vcc));
defparam \D_br_taken_waddr_partial[0] .is_wysiwyg = "true";
defparam \D_br_taken_waddr_partial[0] .power_up = "low";

dffeas D_kill(
	.clk(clk_clk),
	.d(\F_kill~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_kill~q ),
	.prn(vcc));
defparam D_kill.is_wysiwyg = "true";
defparam D_kill.power_up = "low";

cyclonev_lcell_comb \F_ic_tag_rd_addr_nxt[3]~1 (
	.dataa(!\D_issue~q ),
	.datab(!\D_iw_valid~q ),
	.datac(!\D_kill~q ),
	.datad(!\D_ctrl_br~q ),
	.datae(!\D_bht_data[1]~q ),
	.dataf(!\D_ctrl_br_uncond~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_tag_rd_addr_nxt[3]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_tag_rd_addr_nxt[3]~1 .extended_lut = "off";
defparam \F_ic_tag_rd_addr_nxt[3]~1 .lut_mask = 64'hFFFFFDFFFFFFFFFF;
defparam \F_ic_tag_rd_addr_nxt[3]~1 .shared_arith = "off";

cyclonev_lcell_comb \F_ic_data_rd_addr_nxt[0]~0 (
	.dataa(!\D_pc[0]~q ),
	.datab(!\D_br_taken_waddr_partial[0]~q ),
	.datac(!\Add3~1_sumout ),
	.datad(!\D_iw[6]~q ),
	.datae(!\F_ic_tag_rd_addr_nxt[3]~0_combout ),
	.dataf(!\F_ic_tag_rd_addr_nxt[3]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_data_rd_addr_nxt[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_data_rd_addr_nxt[0]~0 .extended_lut = "off";
defparam \F_ic_data_rd_addr_nxt[0]~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \F_ic_data_rd_addr_nxt[0]~0 .shared_arith = "off";

dffeas \E_pc[0] (
	.clk(clk_clk),
	.d(\D_pc[0]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_pc[0]~q ),
	.prn(vcc));
defparam \E_pc[0] .is_wysiwyg = "true";
defparam \E_pc[0] .power_up = "low";

cyclonev_lcell_comb \M_pc_plus_one[0]~0 (
	.dataa(!\E_pc[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_pc_plus_one[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_pc_plus_one[0]~0 .extended_lut = "off";
defparam \M_pc_plus_one[0]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \M_pc_plus_one[0]~0 .shared_arith = "off";

dffeas \M_pc_plus_one[0] (
	.clk(clk_clk),
	.d(\M_pc_plus_one[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_pc_plus_one[0]~q ),
	.prn(vcc));
defparam \M_pc_plus_one[0] .is_wysiwyg = "true";
defparam \M_pc_plus_one[0] .power_up = "low";

dffeas \M_target_pcb[2] (
	.clk(clk_clk),
	.d(\E_src1[2]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_target_pcb[2]~q ),
	.prn(vcc));
defparam \M_target_pcb[2] .is_wysiwyg = "true";
defparam \M_target_pcb[2] .power_up = "low";

dffeas E_ctrl_jmp_indirect(
	.clk(clk_clk),
	.d(\E_ctrl_jmp_indirect_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_ctrl_jmp_indirect~q ),
	.prn(vcc));
defparam E_ctrl_jmp_indirect.is_wysiwyg = "true";
defparam E_ctrl_jmp_indirect.power_up = "low";

dffeas M_ctrl_jmp_indirect(
	.clk(clk_clk),
	.d(\E_ctrl_jmp_indirect~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_ctrl_jmp_indirect~q ),
	.prn(vcc));
defparam M_ctrl_jmp_indirect.is_wysiwyg = "true";
defparam M_ctrl_jmp_indirect.power_up = "low";

cyclonev_lcell_comb \A_pipe_flush_waddr_nxt~0 (
	.dataa(!\M_exc_any~combout ),
	.datab(!\M_pc_plus_one[0]~q ),
	.datac(!\M_target_pcb[2]~q ),
	.datad(!\M_ctrl_jmp_indirect~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_pipe_flush_waddr_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_pipe_flush_waddr_nxt~0 .extended_lut = "off";
defparam \A_pipe_flush_waddr_nxt~0 .lut_mask = 64'hAF3FAF3FAF3FAF3F;
defparam \A_pipe_flush_waddr_nxt~0 .shared_arith = "off";

dffeas \A_pipe_flush_waddr[0] (
	.clk(clk_clk),
	.d(\A_pipe_flush_waddr_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\M_exc_break~0_combout ),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_pipe_flush_waddr[0]~q ),
	.prn(vcc));
defparam \A_pipe_flush_waddr[0] .is_wysiwyg = "true";
defparam \A_pipe_flush_waddr[0] .power_up = "low";

dffeas \D_pc_plus_one[0] (
	.clk(clk_clk),
	.d(\Add3~1_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_pc_plus_one[0]~q ),
	.prn(vcc));
defparam \D_pc_plus_one[0] .is_wysiwyg = "true";
defparam \D_pc_plus_one[0] .power_up = "low";

cyclonev_lcell_comb \E_ctrl_br_cond_nxt~0 (
	.dataa(!\D_iw[4]~q ),
	.datab(!\D_iw[5]~q ),
	.datac(!\D_iw[2]~q ),
	.datad(!\D_iw[3]~q ),
	.datae(!\D_iw[1]~q ),
	.dataf(!\D_iw[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_ctrl_br_cond_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_ctrl_br_cond_nxt~0 .extended_lut = "off";
defparam \E_ctrl_br_cond_nxt~0 .lut_mask = 64'hBFFFFFFF1FFFFFFF;
defparam \E_ctrl_br_cond_nxt~0 .shared_arith = "off";

cyclonev_lcell_comb D_br_pred_not_taken(
	.dataa(!\D_bht_data[1]~q ),
	.datab(!\E_ctrl_br_cond_nxt~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_br_pred_not_taken~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam D_br_pred_not_taken.extended_lut = "off";
defparam D_br_pred_not_taken.lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam D_br_pred_not_taken.shared_arith = "off";

dffeas \E_extra_pc[0] (
	.clk(clk_clk),
	.d(\D_br_taken_waddr_partial[0]~q ),
	.asdata(\D_pc_plus_one[0]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_br_pred_not_taken~combout ),
	.ena(!\A_mem_stall~q ),
	.q(\E_extra_pc[0]~q ),
	.prn(vcc));
defparam \E_extra_pc[0] .is_wysiwyg = "true";
defparam \E_extra_pc[0] .power_up = "low";

dffeas \M_pipe_flush_waddr[0] (
	.clk(clk_clk),
	.d(\E_extra_pc[0]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_pipe_flush_waddr[0]~q ),
	.prn(vcc));
defparam \M_pipe_flush_waddr[0] .is_wysiwyg = "true";
defparam \M_pipe_flush_waddr[0] .power_up = "low";

cyclonev_lcell_comb \F_ic_tag_rd_addr_nxt[3]~2 (
	.dataa(!\A_pipe_flush~q ),
	.datab(!\M_pipe_flush~q ),
	.datac(!\E_valid_jmp_indirect~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_tag_rd_addr_nxt[3]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_tag_rd_addr_nxt[3]~2 .extended_lut = "off";
defparam \F_ic_tag_rd_addr_nxt[3]~2 .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \F_ic_tag_rd_addr_nxt[3]~2 .shared_arith = "off";

cyclonev_lcell_comb \F_ic_tag_rd_addr_nxt[3]~3 (
	.dataa(!\A_pipe_flush~q ),
	.datab(!\M_pipe_flush~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_tag_rd_addr_nxt[3]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_tag_rd_addr_nxt[3]~3 .extended_lut = "off";
defparam \F_ic_tag_rd_addr_nxt[3]~3 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \F_ic_tag_rd_addr_nxt[3]~3 .shared_arith = "off";

cyclonev_lcell_comb \F_ic_data_rd_addr_nxt[0]~1 (
	.dataa(!\F_ic_data_rd_addr_nxt[0]~0_combout ),
	.datab(!\E_src1[2]~q ),
	.datac(!\A_pipe_flush_waddr[0]~q ),
	.datad(!\M_pipe_flush_waddr[0]~q ),
	.datae(!\F_ic_tag_rd_addr_nxt[3]~2_combout ),
	.dataf(!\F_ic_tag_rd_addr_nxt[3]~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_data_rd_addr_nxt[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_data_rd_addr_nxt[0]~1 .extended_lut = "off";
defparam \F_ic_data_rd_addr_nxt[0]~1 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \F_ic_data_rd_addr_nxt[0]~1 .shared_arith = "off";

dffeas \F_pc[0] (
	.clk(clk_clk),
	.d(\F_ic_data_rd_addr_nxt[0]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\F_pc[0]~q ),
	.prn(vcc));
defparam \F_pc[0] .is_wysiwyg = "true";
defparam \F_pc[0] .power_up = "low";

cyclonev_lcell_comb \Add3~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\F_pc[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~5_sumout ),
	.cout(\Add3~6 ),
	.shareout());
defparam \Add3~5 .extended_lut = "off";
defparam \Add3~5 .lut_mask = 64'h00000000000000FF;
defparam \Add3~5 .shared_arith = "off";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[9] ),
	.datae(gnd),
	.dataf(!\Add3~5_sumout ),
	.datag(gnd),
	.cin(\Add0~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~5 .shared_arith = "off";

dffeas \D_br_taken_waddr_partial[1] (
	.clk(clk_clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_br_taken_waddr_partial[1]~q ),
	.prn(vcc));
defparam \D_br_taken_waddr_partial[1] .is_wysiwyg = "true";
defparam \D_br_taken_waddr_partial[1] .power_up = "low";

dffeas \D_iw[7] (
	.clk(clk_clk),
	.d(\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[7] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_iw[7]~q ),
	.prn(vcc));
defparam \D_iw[7] .is_wysiwyg = "true";
defparam \D_iw[7] .power_up = "low";

cyclonev_lcell_comb \F_ic_data_rd_addr_nxt[1]~2 (
	.dataa(!\D_pc[1]~q ),
	.datab(!\D_br_taken_waddr_partial[1]~q ),
	.datac(!\Add3~5_sumout ),
	.datad(!\D_iw[7]~q ),
	.datae(!\F_ic_tag_rd_addr_nxt[3]~0_combout ),
	.dataf(!\F_ic_tag_rd_addr_nxt[3]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_data_rd_addr_nxt[1]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_data_rd_addr_nxt[1]~2 .extended_lut = "off";
defparam \F_ic_data_rd_addr_nxt[1]~2 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \F_ic_data_rd_addr_nxt[1]~2 .shared_arith = "off";

dffeas \E_pc[1] (
	.clk(clk_clk),
	.d(\D_pc[1]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_pc[1]~q ),
	.prn(vcc));
defparam \E_pc[1] .is_wysiwyg = "true";
defparam \E_pc[1] .power_up = "low";

cyclonev_lcell_comb \Add7~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_pc[0]~q ),
	.datae(gnd),
	.dataf(!\E_pc[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add7~1_sumout ),
	.cout(\Add7~2 ),
	.shareout());
defparam \Add7~1 .extended_lut = "off";
defparam \Add7~1 .lut_mask = 64'h0000FF00000000FF;
defparam \Add7~1 .shared_arith = "off";

dffeas \M_pc_plus_one[1] (
	.clk(clk_clk),
	.d(\Add7~1_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_pc_plus_one[1]~q ),
	.prn(vcc));
defparam \M_pc_plus_one[1] .is_wysiwyg = "true";
defparam \M_pc_plus_one[1] .power_up = "low";

dffeas \M_target_pcb[3] (
	.clk(clk_clk),
	.d(\E_src1[3]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_target_pcb[3]~q ),
	.prn(vcc));
defparam \M_target_pcb[3] .is_wysiwyg = "true";
defparam \M_target_pcb[3] .power_up = "low";

cyclonev_lcell_comb \A_pipe_flush_waddr_nxt~1 (
	.dataa(!\M_exc_any~combout ),
	.datab(!\M_pc_plus_one[1]~q ),
	.datac(!\M_ctrl_jmp_indirect~q ),
	.datad(!\M_target_pcb[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_pipe_flush_waddr_nxt~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_pipe_flush_waddr_nxt~1 .extended_lut = "off";
defparam \A_pipe_flush_waddr_nxt~1 .lut_mask = 64'hA3FFA3FFA3FFA3FF;
defparam \A_pipe_flush_waddr_nxt~1 .shared_arith = "off";

dffeas \A_pipe_flush_waddr[1] (
	.clk(clk_clk),
	.d(\A_pipe_flush_waddr_nxt~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\M_exc_break~0_combout ),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_pipe_flush_waddr[1]~q ),
	.prn(vcc));
defparam \A_pipe_flush_waddr[1] .is_wysiwyg = "true";
defparam \A_pipe_flush_waddr[1] .power_up = "low";

dffeas \D_pc_plus_one[1] (
	.clk(clk_clk),
	.d(\Add3~5_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_pc_plus_one[1]~q ),
	.prn(vcc));
defparam \D_pc_plus_one[1] .is_wysiwyg = "true";
defparam \D_pc_plus_one[1] .power_up = "low";

dffeas \E_extra_pc[1] (
	.clk(clk_clk),
	.d(\D_br_taken_waddr_partial[1]~q ),
	.asdata(\D_pc_plus_one[1]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_br_pred_not_taken~combout ),
	.ena(!\A_mem_stall~q ),
	.q(\E_extra_pc[1]~q ),
	.prn(vcc));
defparam \E_extra_pc[1] .is_wysiwyg = "true";
defparam \E_extra_pc[1] .power_up = "low";

dffeas \M_pipe_flush_waddr[1] (
	.clk(clk_clk),
	.d(\E_extra_pc[1]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_pipe_flush_waddr[1]~q ),
	.prn(vcc));
defparam \M_pipe_flush_waddr[1] .is_wysiwyg = "true";
defparam \M_pipe_flush_waddr[1] .power_up = "low";

cyclonev_lcell_comb \F_ic_data_rd_addr_nxt[1]~3 (
	.dataa(!\F_ic_data_rd_addr_nxt[1]~2_combout ),
	.datab(!\E_src1[3]~q ),
	.datac(!\A_pipe_flush_waddr[1]~q ),
	.datad(!\M_pipe_flush_waddr[1]~q ),
	.datae(!\F_ic_tag_rd_addr_nxt[3]~2_combout ),
	.dataf(!\F_ic_tag_rd_addr_nxt[3]~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_data_rd_addr_nxt[1]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_data_rd_addr_nxt[1]~3 .extended_lut = "off";
defparam \F_ic_data_rd_addr_nxt[1]~3 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \F_ic_data_rd_addr_nxt[1]~3 .shared_arith = "off";

dffeas \F_pc[1] (
	.clk(clk_clk),
	.d(\F_ic_data_rd_addr_nxt[1]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\F_pc[1]~q ),
	.prn(vcc));
defparam \F_pc[1] .is_wysiwyg = "true";
defparam \F_pc[1] .power_up = "low";

cyclonev_lcell_comb \Add3~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\F_pc[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~9_sumout ),
	.cout(\Add3~10 ),
	.shareout());
defparam \Add3~9 .extended_lut = "off";
defparam \Add3~9 .lut_mask = 64'h00000000000000FF;
defparam \Add3~9 .shared_arith = "off";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[10] ),
	.datae(gnd),
	.dataf(!\Add3~9_sumout ),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~9 .shared_arith = "off";

dffeas \D_br_taken_waddr_partial[2] (
	.clk(clk_clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_br_taken_waddr_partial[2]~q ),
	.prn(vcc));
defparam \D_br_taken_waddr_partial[2] .is_wysiwyg = "true";
defparam \D_br_taken_waddr_partial[2] .power_up = "low";

dffeas \D_iw[8] (
	.clk(clk_clk),
	.d(\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[8] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_iw[8]~q ),
	.prn(vcc));
defparam \D_iw[8] .is_wysiwyg = "true";
defparam \D_iw[8] .power_up = "low";

cyclonev_lcell_comb \F_ic_data_rd_addr_nxt[2]~4 (
	.dataa(!\D_pc[2]~q ),
	.datab(!\D_br_taken_waddr_partial[2]~q ),
	.datac(!\Add3~9_sumout ),
	.datad(!\D_iw[8]~q ),
	.datae(!\F_ic_tag_rd_addr_nxt[3]~0_combout ),
	.dataf(!\F_ic_tag_rd_addr_nxt[3]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_data_rd_addr_nxt[2]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_data_rd_addr_nxt[2]~4 .extended_lut = "off";
defparam \F_ic_data_rd_addr_nxt[2]~4 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \F_ic_data_rd_addr_nxt[2]~4 .shared_arith = "off";

dffeas \E_pc[2] (
	.clk(clk_clk),
	.d(\D_pc[2]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_pc[2]~q ),
	.prn(vcc));
defparam \E_pc[2] .is_wysiwyg = "true";
defparam \E_pc[2] .power_up = "low";

cyclonev_lcell_comb \Add7~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_pc[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add7~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add7~5_sumout ),
	.cout(\Add7~6 ),
	.shareout());
defparam \Add7~5 .extended_lut = "off";
defparam \Add7~5 .lut_mask = 64'h00000000000000FF;
defparam \Add7~5 .shared_arith = "off";

dffeas \M_pc_plus_one[2] (
	.clk(clk_clk),
	.d(\Add7~5_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_pc_plus_one[2]~q ),
	.prn(vcc));
defparam \M_pc_plus_one[2] .is_wysiwyg = "true";
defparam \M_pc_plus_one[2] .power_up = "low";

dffeas \M_target_pcb[4] (
	.clk(clk_clk),
	.d(\E_src1[4]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_target_pcb[4]~q ),
	.prn(vcc));
defparam \M_target_pcb[4] .is_wysiwyg = "true";
defparam \M_target_pcb[4] .power_up = "low";

cyclonev_lcell_comb \A_pipe_flush_waddr_nxt~2 (
	.dataa(!\M_exc_any~combout ),
	.datab(!\M_pc_plus_one[2]~q ),
	.datac(!\M_ctrl_jmp_indirect~q ),
	.datad(!\M_target_pcb[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_pipe_flush_waddr_nxt~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_pipe_flush_waddr_nxt~2 .extended_lut = "off";
defparam \A_pipe_flush_waddr_nxt~2 .lut_mask = 64'hA3FFA3FFA3FFA3FF;
defparam \A_pipe_flush_waddr_nxt~2 .shared_arith = "off";

dffeas \A_pipe_flush_waddr[2] (
	.clk(clk_clk),
	.d(\A_pipe_flush_waddr_nxt~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\M_exc_break~0_combout ),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_pipe_flush_waddr[2]~q ),
	.prn(vcc));
defparam \A_pipe_flush_waddr[2] .is_wysiwyg = "true";
defparam \A_pipe_flush_waddr[2] .power_up = "low";

dffeas \D_pc_plus_one[2] (
	.clk(clk_clk),
	.d(\Add3~9_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_pc_plus_one[2]~q ),
	.prn(vcc));
defparam \D_pc_plus_one[2] .is_wysiwyg = "true";
defparam \D_pc_plus_one[2] .power_up = "low";

dffeas \E_extra_pc[2] (
	.clk(clk_clk),
	.d(\D_br_taken_waddr_partial[2]~q ),
	.asdata(\D_pc_plus_one[2]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_br_pred_not_taken~combout ),
	.ena(!\A_mem_stall~q ),
	.q(\E_extra_pc[2]~q ),
	.prn(vcc));
defparam \E_extra_pc[2] .is_wysiwyg = "true";
defparam \E_extra_pc[2] .power_up = "low";

dffeas \M_pipe_flush_waddr[2] (
	.clk(clk_clk),
	.d(\E_extra_pc[2]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_pipe_flush_waddr[2]~q ),
	.prn(vcc));
defparam \M_pipe_flush_waddr[2] .is_wysiwyg = "true";
defparam \M_pipe_flush_waddr[2] .power_up = "low";

cyclonev_lcell_comb \F_ic_data_rd_addr_nxt[2]~5 (
	.dataa(!\F_ic_data_rd_addr_nxt[2]~4_combout ),
	.datab(!\E_src1[4]~q ),
	.datac(!\A_pipe_flush_waddr[2]~q ),
	.datad(!\M_pipe_flush_waddr[2]~q ),
	.datae(!\F_ic_tag_rd_addr_nxt[3]~2_combout ),
	.dataf(!\F_ic_tag_rd_addr_nxt[3]~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_data_rd_addr_nxt[2]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_data_rd_addr_nxt[2]~5 .extended_lut = "off";
defparam \F_ic_data_rd_addr_nxt[2]~5 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \F_ic_data_rd_addr_nxt[2]~5 .shared_arith = "off";

dffeas \F_pc[2] (
	.clk(clk_clk),
	.d(\F_ic_data_rd_addr_nxt[2]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\F_pc[2]~q ),
	.prn(vcc));
defparam \F_pc[2] .is_wysiwyg = "true";
defparam \F_pc[2] .power_up = "low";

cyclonev_lcell_comb \F_ic_valid~4 (
	.dataa(!\first_nios2_system_cpu_cpu_ic_tag|the_altsyncram|auto_generated|q_b[7] ),
	.datab(!\first_nios2_system_cpu_cpu_ic_tag|the_altsyncram|auto_generated|q_b[9] ),
	.datac(!\first_nios2_system_cpu_cpu_ic_tag|the_altsyncram|auto_generated|q_b[8] ),
	.datad(!\F_pc[0]~q ),
	.datae(!\F_pc[1]~q ),
	.dataf(!\F_pc[2]~q ),
	.datag(!\first_nios2_system_cpu_cpu_ic_tag|the_altsyncram|auto_generated|q_b[6] ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_valid~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_valid~4 .extended_lut = "on";
defparam \F_ic_valid~4 .lut_mask = 64'hFAFCFAFCFAFCFAFC;
defparam \F_ic_valid~4 .shared_arith = "off";

cyclonev_lcell_comb \F_ic_valid~0 (
	.dataa(!\first_nios2_system_cpu_cpu_ic_tag|the_altsyncram|auto_generated|q_b[11] ),
	.datab(!\first_nios2_system_cpu_cpu_ic_tag|the_altsyncram|auto_generated|q_b[13] ),
	.datac(!\first_nios2_system_cpu_cpu_ic_tag|the_altsyncram|auto_generated|q_b[12] ),
	.datad(!\F_pc[2]~q ),
	.datae(!\F_pc[1]~q ),
	.dataf(!\F_ic_valid~4_combout ),
	.datag(!\first_nios2_system_cpu_cpu_ic_tag|the_altsyncram|auto_generated|q_b[10] ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_valid~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_valid~0 .extended_lut = "on";
defparam \F_ic_valid~0 .lut_mask = 64'hFAFCFAFCFAFCFAFC;
defparam \F_ic_valid~0 .shared_arith = "off";

dffeas \D_pc[14] (
	.clk(clk_clk),
	.d(\F_pc[14]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_pc[14]~q ),
	.prn(vcc));
defparam \D_pc[14] .is_wysiwyg = "true";
defparam \D_pc[14] .power_up = "low";

dffeas \D_pc[13] (
	.clk(clk_clk),
	.d(\F_pc[13]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_pc[13]~q ),
	.prn(vcc));
defparam \D_pc[13] .is_wysiwyg = "true";
defparam \D_pc[13] .power_up = "low";

dffeas \D_pc[12] (
	.clk(clk_clk),
	.d(\F_pc[12]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_pc[12]~q ),
	.prn(vcc));
defparam \D_pc[12] .is_wysiwyg = "true";
defparam \D_pc[12] .power_up = "low";

dffeas \D_pc[11] (
	.clk(clk_clk),
	.d(\F_pc[11]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_pc[11]~q ),
	.prn(vcc));
defparam \D_pc[11] .is_wysiwyg = "true";
defparam \D_pc[11] .power_up = "low";

dffeas \D_pc[10] (
	.clk(clk_clk),
	.d(\F_pc[10]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_pc[10]~q ),
	.prn(vcc));
defparam \D_pc[10] .is_wysiwyg = "true";
defparam \D_pc[10] .power_up = "low";

dffeas \D_pc[9] (
	.clk(clk_clk),
	.d(\F_pc[9]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_pc[9]~q ),
	.prn(vcc));
defparam \D_pc[9] .is_wysiwyg = "true";
defparam \D_pc[9] .power_up = "low";

dffeas \D_pc[8] (
	.clk(clk_clk),
	.d(\F_pc[8]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_pc[8]~q ),
	.prn(vcc));
defparam \D_pc[8] .is_wysiwyg = "true";
defparam \D_pc[8] .power_up = "low";

dffeas \D_pc[7] (
	.clk(clk_clk),
	.d(\F_pc[7]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_pc[7]~q ),
	.prn(vcc));
defparam \D_pc[7] .is_wysiwyg = "true";
defparam \D_pc[7] .power_up = "low";

dffeas \D_pc[6] (
	.clk(clk_clk),
	.d(\F_pc[6]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_pc[6]~q ),
	.prn(vcc));
defparam \D_pc[6] .is_wysiwyg = "true";
defparam \D_pc[6] .power_up = "low";

dffeas \D_pc[5] (
	.clk(clk_clk),
	.d(\F_pc[5]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_pc[5]~q ),
	.prn(vcc));
defparam \D_pc[5] .is_wysiwyg = "true";
defparam \D_pc[5] .power_up = "low";

dffeas \D_pc[4] (
	.clk(clk_clk),
	.d(\F_pc[4]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_pc[4]~q ),
	.prn(vcc));
defparam \D_pc[4] .is_wysiwyg = "true";
defparam \D_pc[4] .power_up = "low";

cyclonev_lcell_comb \Add3~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\F_pc[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~13_sumout ),
	.cout(\Add3~14 ),
	.shareout());
defparam \Add3~13 .extended_lut = "off";
defparam \Add3~13 .lut_mask = 64'h00000000000000FF;
defparam \Add3~13 .shared_arith = "off";

cyclonev_lcell_comb \Add3~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\F_pc[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~17_sumout ),
	.cout(\Add3~18 ),
	.shareout());
defparam \Add3~17 .extended_lut = "off";
defparam \Add3~17 .lut_mask = 64'h00000000000000FF;
defparam \Add3~17 .shared_arith = "off";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[11] ),
	.datae(gnd),
	.dataf(!\Add3~13_sumout ),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~13 .shared_arith = "off";

cyclonev_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[12] ),
	.datae(gnd),
	.dataf(!\Add3~17_sumout ),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~17 .shared_arith = "off";

dffeas \D_br_taken_waddr_partial[4] (
	.clk(clk_clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_br_taken_waddr_partial[4]~q ),
	.prn(vcc));
defparam \D_br_taken_waddr_partial[4] .is_wysiwyg = "true";
defparam \D_br_taken_waddr_partial[4] .power_up = "low";

dffeas \D_iw[10] (
	.clk(clk_clk),
	.d(\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[10] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_iw[10]~q ),
	.prn(vcc));
defparam \D_iw[10] .is_wysiwyg = "true";
defparam \D_iw[10] .power_up = "low";

cyclonev_lcell_comb \F_ic_tag_rd_addr_nxt[1]~6 (
	.dataa(!\D_pc[4]~q ),
	.datab(!\D_br_taken_waddr_partial[4]~q ),
	.datac(!\Add3~17_sumout ),
	.datad(!\D_iw[10]~q ),
	.datae(!\F_ic_tag_rd_addr_nxt[3]~0_combout ),
	.dataf(!\F_ic_tag_rd_addr_nxt[3]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_tag_rd_addr_nxt[1]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_tag_rd_addr_nxt[1]~6 .extended_lut = "off";
defparam \F_ic_tag_rd_addr_nxt[1]~6 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \F_ic_tag_rd_addr_nxt[1]~6 .shared_arith = "off";

dffeas \E_pc[4] (
	.clk(clk_clk),
	.d(\D_pc[4]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_pc[4]~q ),
	.prn(vcc));
defparam \E_pc[4] .is_wysiwyg = "true";
defparam \E_pc[4] .power_up = "low";

dffeas \E_pc[3] (
	.clk(clk_clk),
	.d(\D_pc[3]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_pc[3]~q ),
	.prn(vcc));
defparam \E_pc[3] .is_wysiwyg = "true";
defparam \E_pc[3] .power_up = "low";

cyclonev_lcell_comb \Add7~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_pc[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add7~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add7~9_sumout ),
	.cout(\Add7~10 ),
	.shareout());
defparam \Add7~9 .extended_lut = "off";
defparam \Add7~9 .lut_mask = 64'h00000000000000FF;
defparam \Add7~9 .shared_arith = "off";

cyclonev_lcell_comb \Add7~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_pc[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add7~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add7~13_sumout ),
	.cout(\Add7~14 ),
	.shareout());
defparam \Add7~13 .extended_lut = "off";
defparam \Add7~13 .lut_mask = 64'h00000000000000FF;
defparam \Add7~13 .shared_arith = "off";

dffeas \M_pc_plus_one[4] (
	.clk(clk_clk),
	.d(\Add7~13_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_pc_plus_one[4]~q ),
	.prn(vcc));
defparam \M_pc_plus_one[4] .is_wysiwyg = "true";
defparam \M_pc_plus_one[4] .power_up = "low";

dffeas \M_target_pcb[6] (
	.clk(clk_clk),
	.d(\E_src1[6]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_target_pcb[6]~q ),
	.prn(vcc));
defparam \M_target_pcb[6] .is_wysiwyg = "true";
defparam \M_target_pcb[6] .power_up = "low";

cyclonev_lcell_comb \A_pipe_flush_waddr_nxt~4 (
	.dataa(!\M_exc_any~combout ),
	.datab(!\M_pc_plus_one[4]~q ),
	.datac(!\M_ctrl_jmp_indirect~q ),
	.datad(!\M_target_pcb[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_pipe_flush_waddr_nxt~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_pipe_flush_waddr_nxt~4 .extended_lut = "off";
defparam \A_pipe_flush_waddr_nxt~4 .lut_mask = 64'hA3FFA3FFA3FFA3FF;
defparam \A_pipe_flush_waddr_nxt~4 .shared_arith = "off";

dffeas \A_pipe_flush_waddr[4] (
	.clk(clk_clk),
	.d(\A_pipe_flush_waddr_nxt~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\M_exc_break~0_combout ),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_pipe_flush_waddr[4]~q ),
	.prn(vcc));
defparam \A_pipe_flush_waddr[4] .is_wysiwyg = "true";
defparam \A_pipe_flush_waddr[4] .power_up = "low";

dffeas \D_pc_plus_one[4] (
	.clk(clk_clk),
	.d(\Add3~17_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_pc_plus_one[4]~q ),
	.prn(vcc));
defparam \D_pc_plus_one[4] .is_wysiwyg = "true";
defparam \D_pc_plus_one[4] .power_up = "low";

dffeas \E_extra_pc[4] (
	.clk(clk_clk),
	.d(\D_br_taken_waddr_partial[4]~q ),
	.asdata(\D_pc_plus_one[4]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_br_pred_not_taken~combout ),
	.ena(!\A_mem_stall~q ),
	.q(\E_extra_pc[4]~q ),
	.prn(vcc));
defparam \E_extra_pc[4] .is_wysiwyg = "true";
defparam \E_extra_pc[4] .power_up = "low";

dffeas \M_pipe_flush_waddr[4] (
	.clk(clk_clk),
	.d(\E_extra_pc[4]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_pipe_flush_waddr[4]~q ),
	.prn(vcc));
defparam \M_pipe_flush_waddr[4] .is_wysiwyg = "true";
defparam \M_pipe_flush_waddr[4] .power_up = "low";

cyclonev_lcell_comb \F_ic_tag_rd_addr_nxt[1]~7 (
	.dataa(!\F_ic_tag_rd_addr_nxt[1]~6_combout ),
	.datab(!\E_src1[6]~q ),
	.datac(!\A_pipe_flush_waddr[4]~q ),
	.datad(!\M_pipe_flush_waddr[4]~q ),
	.datae(!\F_ic_tag_rd_addr_nxt[3]~2_combout ),
	.dataf(!\F_ic_tag_rd_addr_nxt[3]~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_tag_rd_addr_nxt[1]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_tag_rd_addr_nxt[1]~7 .extended_lut = "off";
defparam \F_ic_tag_rd_addr_nxt[1]~7 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \F_ic_tag_rd_addr_nxt[1]~7 .shared_arith = "off";

dffeas \F_pc[4] (
	.clk(clk_clk),
	.d(\F_ic_tag_rd_addr_nxt[1]~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\F_pc[4]~q ),
	.prn(vcc));
defparam \F_pc[4] .is_wysiwyg = "true";
defparam \F_pc[4] .power_up = "low";

cyclonev_lcell_comb \Add3~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\F_pc[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~21_sumout ),
	.cout(\Add3~22 ),
	.shareout());
defparam \Add3~21 .extended_lut = "off";
defparam \Add3~21 .lut_mask = 64'h00000000000000FF;
defparam \Add3~21 .shared_arith = "off";

cyclonev_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[13] ),
	.datae(gnd),
	.dataf(!\Add3~21_sumout ),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~21 .shared_arith = "off";

dffeas \D_br_taken_waddr_partial[5] (
	.clk(clk_clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_br_taken_waddr_partial[5]~q ),
	.prn(vcc));
defparam \D_br_taken_waddr_partial[5] .is_wysiwyg = "true";
defparam \D_br_taken_waddr_partial[5] .power_up = "low";

cyclonev_lcell_comb \F_ic_tag_rd_addr_nxt[2]~8 (
	.dataa(!\D_pc[5]~q ),
	.datab(!\D_br_taken_waddr_partial[5]~q ),
	.datac(!\Add3~21_sumout ),
	.datad(!\D_iw[11]~q ),
	.datae(!\F_ic_tag_rd_addr_nxt[3]~0_combout ),
	.dataf(!\F_ic_tag_rd_addr_nxt[3]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_tag_rd_addr_nxt[2]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_tag_rd_addr_nxt[2]~8 .extended_lut = "off";
defparam \F_ic_tag_rd_addr_nxt[2]~8 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \F_ic_tag_rd_addr_nxt[2]~8 .shared_arith = "off";

dffeas \E_pc[5] (
	.clk(clk_clk),
	.d(\D_pc[5]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_pc[5]~q ),
	.prn(vcc));
defparam \E_pc[5] .is_wysiwyg = "true";
defparam \E_pc[5] .power_up = "low";

cyclonev_lcell_comb \Add7~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_pc[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add7~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add7~17_sumout ),
	.cout(\Add7~18 ),
	.shareout());
defparam \Add7~17 .extended_lut = "off";
defparam \Add7~17 .lut_mask = 64'h00000000000000FF;
defparam \Add7~17 .shared_arith = "off";

dffeas \M_pc_plus_one[5] (
	.clk(clk_clk),
	.d(\Add7~17_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_pc_plus_one[5]~q ),
	.prn(vcc));
defparam \M_pc_plus_one[5] .is_wysiwyg = "true";
defparam \M_pc_plus_one[5] .power_up = "low";

dffeas \M_target_pcb[7] (
	.clk(clk_clk),
	.d(\E_src1[7]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_target_pcb[7]~q ),
	.prn(vcc));
defparam \M_target_pcb[7] .is_wysiwyg = "true";
defparam \M_target_pcb[7] .power_up = "low";

cyclonev_lcell_comb \A_pipe_flush_waddr_nxt~5 (
	.dataa(!\M_exc_any~combout ),
	.datab(!\M_pc_plus_one[5]~q ),
	.datac(!\M_ctrl_jmp_indirect~q ),
	.datad(!\M_target_pcb[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_pipe_flush_waddr_nxt~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_pipe_flush_waddr_nxt~5 .extended_lut = "off";
defparam \A_pipe_flush_waddr_nxt~5 .lut_mask = 64'hA3FFA3FFA3FFA3FF;
defparam \A_pipe_flush_waddr_nxt~5 .shared_arith = "off";

dffeas \A_pipe_flush_waddr[5] (
	.clk(clk_clk),
	.d(\A_pipe_flush_waddr_nxt~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\M_exc_break~0_combout ),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_pipe_flush_waddr[5]~q ),
	.prn(vcc));
defparam \A_pipe_flush_waddr[5] .is_wysiwyg = "true";
defparam \A_pipe_flush_waddr[5] .power_up = "low";

dffeas \D_pc_plus_one[5] (
	.clk(clk_clk),
	.d(\Add3~21_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_pc_plus_one[5]~q ),
	.prn(vcc));
defparam \D_pc_plus_one[5] .is_wysiwyg = "true";
defparam \D_pc_plus_one[5] .power_up = "low";

dffeas \E_extra_pc[5] (
	.clk(clk_clk),
	.d(\D_br_taken_waddr_partial[5]~q ),
	.asdata(\D_pc_plus_one[5]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_br_pred_not_taken~combout ),
	.ena(!\A_mem_stall~q ),
	.q(\E_extra_pc[5]~q ),
	.prn(vcc));
defparam \E_extra_pc[5] .is_wysiwyg = "true";
defparam \E_extra_pc[5] .power_up = "low";

dffeas \M_pipe_flush_waddr[5] (
	.clk(clk_clk),
	.d(\E_extra_pc[5]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_pipe_flush_waddr[5]~q ),
	.prn(vcc));
defparam \M_pipe_flush_waddr[5] .is_wysiwyg = "true";
defparam \M_pipe_flush_waddr[5] .power_up = "low";

cyclonev_lcell_comb \F_ic_tag_rd_addr_nxt[2]~9 (
	.dataa(!\F_ic_tag_rd_addr_nxt[2]~8_combout ),
	.datab(!\E_src1[7]~q ),
	.datac(!\A_pipe_flush_waddr[5]~q ),
	.datad(!\M_pipe_flush_waddr[5]~q ),
	.datae(!\F_ic_tag_rd_addr_nxt[3]~2_combout ),
	.dataf(!\F_ic_tag_rd_addr_nxt[3]~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_tag_rd_addr_nxt[2]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_tag_rd_addr_nxt[2]~9 .extended_lut = "off";
defparam \F_ic_tag_rd_addr_nxt[2]~9 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \F_ic_tag_rd_addr_nxt[2]~9 .shared_arith = "off";

dffeas \F_pc[5] (
	.clk(clk_clk),
	.d(\F_ic_tag_rd_addr_nxt[2]~9_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\F_pc[5]~q ),
	.prn(vcc));
defparam \F_pc[5] .is_wysiwyg = "true";
defparam \F_pc[5] .power_up = "low";

cyclonev_lcell_comb \Add3~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\F_pc[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~25_sumout ),
	.cout(\Add3~26 ),
	.shareout());
defparam \Add3~25 .extended_lut = "off";
defparam \Add3~25 .lut_mask = 64'h00000000000000FF;
defparam \Add3~25 .shared_arith = "off";

cyclonev_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[14] ),
	.datae(gnd),
	.dataf(!\Add3~25_sumout ),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout());
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~33 .shared_arith = "off";

dffeas \D_br_taken_waddr_partial[6] (
	.clk(clk_clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_br_taken_waddr_partial[6]~q ),
	.prn(vcc));
defparam \D_br_taken_waddr_partial[6] .is_wysiwyg = "true";
defparam \D_br_taken_waddr_partial[6] .power_up = "low";

cyclonev_lcell_comb \F_ic_tag_rd_addr_nxt[3]~10 (
	.dataa(!\D_pc[6]~q ),
	.datab(!\D_br_taken_waddr_partial[6]~q ),
	.datac(!\Add3~25_sumout ),
	.datad(!\D_iw[12]~q ),
	.datae(!\F_ic_tag_rd_addr_nxt[3]~0_combout ),
	.dataf(!\F_ic_tag_rd_addr_nxt[3]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_tag_rd_addr_nxt[3]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_tag_rd_addr_nxt[3]~10 .extended_lut = "off";
defparam \F_ic_tag_rd_addr_nxt[3]~10 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \F_ic_tag_rd_addr_nxt[3]~10 .shared_arith = "off";

cyclonev_lcell_comb \A_slow_inst_result_nxt[8]~40 (
	.dataa(!\d_readdata_d1[8]~q ),
	.datab(!\d_readdata_d1[24]~q ),
	.datac(!\A_slow_inst_result[9]~0_combout ),
	.datad(!\A_slow_inst_result[9]~1_combout ),
	.datae(!src0_valid),
	.dataf(!av_readdata_pre_8),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[8]~40_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[8]~40 .extended_lut = "off";
defparam \A_slow_inst_result_nxt[8]~40 .lut_mask = 64'h7FF7FFFFFFFFFFFF;
defparam \A_slow_inst_result_nxt[8]~40 .shared_arith = "off";

cyclonev_lcell_comb \A_slow_inst_result_nxt[8]~68 (
	.dataa(!\A_slow_inst_result_nxt[8]~40_combout ),
	.datab(!q_a_8),
	.datac(!\A_slow_ld_data_fill_bit~0_combout ),
	.datad(!src0_valid1),
	.datae(!\A_slow_inst_result[9]~0_combout ),
	.dataf(!\A_slow_inst_result[9]~1_combout ),
	.datag(!src_payload7),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[8]~68_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[8]~68 .extended_lut = "on";
defparam \A_slow_inst_result_nxt[8]~68 .lut_mask = 64'hFFD8FFD8FFD8FFD8;
defparam \A_slow_inst_result_nxt[8]~68 .shared_arith = "off";

dffeas \A_slow_inst_result[8] (
	.clk(clk_clk),
	.d(\A_slow_inst_result_nxt[8]~68_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_ctrl_ld~q ),
	.q(\A_slow_inst_result[8]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[8] .is_wysiwyg = "true";
defparam \A_slow_inst_result[8] .power_up = "low";

cyclonev_lcell_comb \E_rot_mask[0]~0 (
	.dataa(!\E_src2[2]~q ),
	.datab(!\E_src2[1]~q ),
	.datac(!\E_src2[0]~q ),
	.datad(!\E_ctrl_shift_rot_right~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_mask[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_mask[0]~0 .extended_lut = "off";
defparam \E_rot_mask[0]~0 .lut_mask = 64'hFF7FFF7FFF7FFF7F;
defparam \E_rot_mask[0]~0 .shared_arith = "off";

dffeas \M_rot_mask[0] (
	.clk(clk_clk),
	.d(\E_rot_mask[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_rot_mask[0]~q ),
	.prn(vcc));
defparam \M_rot_mask[0] .is_wysiwyg = "true";
defparam \M_rot_mask[0] .power_up = "low";

cyclonev_lcell_comb \E_rot_step1[4]~6 (
	.dataa(!\E_src1[4]~q ),
	.datab(!\E_src1[3]~q ),
	.datac(!\E_src1[2]~q ),
	.datad(!\E_src1[1]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add10~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[4]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[4]~6 .extended_lut = "off";
defparam \E_rot_step1[4]~6 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[4]~6 .shared_arith = "off";

cyclonev_lcell_comb \E_rot_step1[8]~7 (
	.dataa(!\E_src1[8]~q ),
	.datab(!\E_src1[7]~q ),
	.datac(!\E_src1[6]~q ),
	.datad(!\E_src1[5]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add10~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[8]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[8]~7 .extended_lut = "off";
defparam \E_rot_step1[8]~7 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[8]~7 .shared_arith = "off";

cyclonev_lcell_comb \Add10~1 (
	.dataa(!\E_src2[2]~q ),
	.datab(!\E_src2[1]~q ),
	.datac(!\E_src2[0]~q ),
	.datad(!\E_ctrl_shift_rot_right~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add10~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add10~1 .extended_lut = "off";
defparam \Add10~1 .lut_mask = 64'h6996699669966996;
defparam \Add10~1 .shared_arith = "off";

dffeas \M_rot_prestep2[8] (
	.clk(clk_clk),
	.d(\E_rot_step1[4]~6_combout ),
	.asdata(\E_rot_step1[8]~7_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add10~1_combout ),
	.ena(!\A_mem_stall~q ),
	.q(\M_rot_prestep2[8]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[8] .is_wysiwyg = "true";
defparam \M_rot_prestep2[8] .power_up = "low";

cyclonev_lcell_comb \E_rot_step1[28]~0 (
	.dataa(!\E_src1[28]~q ),
	.datab(!\E_src1[27]~q ),
	.datac(!\E_src1[26]~q ),
	.datad(!\E_src1[25]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add10~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[28]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[28]~0 .extended_lut = "off";
defparam \E_rot_step1[28]~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[28]~0 .shared_arith = "off";

cyclonev_lcell_comb \E_rot_step1[0]~1 (
	.dataa(!\E_src1[0]~q ),
	.datab(!\E_src1[31]~q ),
	.datac(!\E_src1[30]~q ),
	.datad(!\E_src1[29]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add10~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[0]~1 .extended_lut = "off";
defparam \E_rot_step1[0]~1 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[0]~1 .shared_arith = "off";

dffeas \M_rot_prestep2[0] (
	.clk(clk_clk),
	.d(\E_rot_step1[28]~0_combout ),
	.asdata(\E_rot_step1[0]~1_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add10~1_combout ),
	.ena(!\A_mem_stall~q ),
	.q(\M_rot_prestep2[0]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[0] .is_wysiwyg = "true";
defparam \M_rot_prestep2[0] .power_up = "low";

cyclonev_lcell_comb \A_slow_inst_result_nxt[20]~34 (
	.dataa(!\A_ctrl_ld32~q ),
	.datab(!\d_readdata_d1[20]~q ),
	.datac(!read_latency_shift_reg_01),
	.datad(!src0_valid),
	.datae(!av_readdata_pre_20),
	.dataf(!av_readdata_pre_201),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[20]~34_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[20]~34 .extended_lut = "off";
defparam \A_slow_inst_result_nxt[20]~34 .lut_mask = 64'h27FFFFFFFFFFFFFF;
defparam \A_slow_inst_result_nxt[20]~34 .shared_arith = "off";

cyclonev_lcell_comb \A_slow_inst_result_nxt[20]~17 (
	.dataa(!\A_ctrl_ld32~q ),
	.datab(!\A_ld_align_byte2_byte3_fill~q ),
	.datac(!\A_slow_ld_data_fill_bit~0_combout ),
	.datad(!src0_valid1),
	.datae(!q_a_20),
	.dataf(!\A_slow_inst_result_nxt[20]~34_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[20]~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[20]~17 .extended_lut = "off";
defparam \A_slow_inst_result_nxt[20]~17 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \A_slow_inst_result_nxt[20]~17 .shared_arith = "off";

dffeas \A_slow_inst_result[20] (
	.clk(clk_clk),
	.d(\A_slow_inst_result_nxt[20]~17_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_ctrl_ld~q ),
	.q(\A_slow_inst_result[20]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[20] .is_wysiwyg = "true";
defparam \A_slow_inst_result[20] .power_up = "low";

cyclonev_lcell_comb \A_slow_inst_result_nxt[16]~29 (
	.dataa(!\A_ctrl_ld32~q ),
	.datab(!\A_ld_align_byte2_byte3_fill~q ),
	.datac(!src0_valid),
	.datad(!av_readdata_pre_16),
	.datae(!src_payload11),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[16]~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[16]~29 .extended_lut = "off";
defparam \A_slow_inst_result_nxt[16]~29 .lut_mask = 64'hFFD8FFFFFFD8FFFF;
defparam \A_slow_inst_result_nxt[16]~29 .shared_arith = "off";

cyclonev_lcell_comb \A_slow_inst_result_nxt[16]~22 (
	.dataa(!\A_ctrl_ld32~q ),
	.datab(!\d_readdata_d1[16]~q ),
	.datac(!\A_slow_ld_data_fill_bit~0_combout ),
	.datad(!src0_valid1),
	.datae(!q_a_16),
	.dataf(!\A_slow_inst_result_nxt[16]~29_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[16]~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[16]~22 .extended_lut = "off";
defparam \A_slow_inst_result_nxt[16]~22 .lut_mask = 64'h7FFFFFFFBFFFFFFF;
defparam \A_slow_inst_result_nxt[16]~22 .shared_arith = "off";

dffeas \A_slow_inst_result[16] (
	.clk(clk_clk),
	.d(\A_slow_inst_result_nxt[16]~22_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_ctrl_ld~q ),
	.q(\A_slow_inst_result[16]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[16] .is_wysiwyg = "true";
defparam \A_slow_inst_result[16] .power_up = "low";

cyclonev_lcell_comb \A_slow_inst_result_nxt[12]~44 (
	.dataa(!\d_readdata_d1[12]~q ),
	.datab(!\d_readdata_d1[28]~q ),
	.datac(!\A_slow_inst_result[9]~0_combout ),
	.datad(!\A_slow_inst_result[9]~1_combout ),
	.datae(!src0_valid),
	.dataf(!av_readdata_pre_12),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[12]~44_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[12]~44 .extended_lut = "off";
defparam \A_slow_inst_result_nxt[12]~44 .lut_mask = 64'h7FF7FFFFFFFFFFFF;
defparam \A_slow_inst_result_nxt[12]~44 .shared_arith = "off";

cyclonev_lcell_comb \A_slow_inst_result_nxt[12]~56 (
	.dataa(!\A_slow_inst_result[9]~1_combout ),
	.datab(!\A_slow_inst_result_nxt[12]~44_combout ),
	.datac(!\A_slow_ld_data_fill_bit~0_combout ),
	.datad(!src_payload13),
	.datae(!\A_slow_inst_result[9]~0_combout ),
	.dataf(!q_a_12),
	.datag(!src0_valid1),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[12]~56_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[12]~56 .extended_lut = "on";
defparam \A_slow_inst_result_nxt[12]~56 .lut_mask = 64'hFFD8FFD8FFD8FFD8;
defparam \A_slow_inst_result_nxt[12]~56 .shared_arith = "off";

dffeas \A_slow_inst_result[12] (
	.clk(clk_clk),
	.d(\A_slow_inst_result_nxt[12]~56_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_ctrl_ld~q ),
	.q(\A_slow_inst_result[12]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[12] .is_wysiwyg = "true";
defparam \A_slow_inst_result[12] .power_up = "low";

dffeas \M_rot_prestep2[12] (
	.clk(clk_clk),
	.d(\E_rot_step1[8]~7_combout ),
	.asdata(\E_rot_step1[12]~4_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add10~1_combout ),
	.ena(!\A_mem_stall~q ),
	.q(\M_rot_prestep2[12]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[12] .is_wysiwyg = "true";
defparam \M_rot_prestep2[12] .power_up = "low";

dffeas \M_rot_prestep2[4] (
	.clk(clk_clk),
	.d(\E_rot_step1[0]~1_combout ),
	.asdata(\E_rot_step1[4]~6_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add10~1_combout ),
	.ena(!\A_mem_stall~q ),
	.q(\M_rot_prestep2[4]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[4] .is_wysiwyg = "true";
defparam \M_rot_prestep2[4] .power_up = "low";

cyclonev_lcell_comb \A_slow_inst_result_nxt[21]~27 (
	.dataa(!\A_ctrl_ld32~q ),
	.datab(!\A_ld_align_byte2_byte3_fill~q ),
	.datac(!src0_valid),
	.datad(!av_readdata_pre_21),
	.datae(!src_payload4),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[21]~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[21]~27 .extended_lut = "off";
defparam \A_slow_inst_result_nxt[21]~27 .lut_mask = 64'hFFD8FFFFFFD8FFFF;
defparam \A_slow_inst_result_nxt[21]~27 .shared_arith = "off";

cyclonev_lcell_comb \A_slow_inst_result_nxt[21]~13 (
	.dataa(!\A_ctrl_ld32~q ),
	.datab(!\d_readdata_d1[21]~q ),
	.datac(!\A_slow_ld_data_fill_bit~0_combout ),
	.datad(!src0_valid1),
	.datae(!q_a_21),
	.dataf(!\A_slow_inst_result_nxt[21]~27_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[21]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[21]~13 .extended_lut = "off";
defparam \A_slow_inst_result_nxt[21]~13 .lut_mask = 64'h7FFFFFFFBFFFFFFF;
defparam \A_slow_inst_result_nxt[21]~13 .shared_arith = "off";

dffeas \A_slow_inst_result[21] (
	.clk(clk_clk),
	.d(\A_slow_inst_result_nxt[21]~13_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_ctrl_ld~q ),
	.q(\A_slow_inst_result[21]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[21] .is_wysiwyg = "true";
defparam \A_slow_inst_result[21] .power_up = "low";

cyclonev_lcell_comb \A_slow_inst_result_nxt[17]~30 (
	.dataa(!\A_ctrl_ld32~q ),
	.datab(!\A_ld_align_byte2_byte3_fill~q ),
	.datac(!src0_valid),
	.datad(!av_readdata_pre_17),
	.datae(!src_payload9),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[17]~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[17]~30 .extended_lut = "off";
defparam \A_slow_inst_result_nxt[17]~30 .lut_mask = 64'hFFD8FFFFFFD8FFFF;
defparam \A_slow_inst_result_nxt[17]~30 .shared_arith = "off";

cyclonev_lcell_comb \A_slow_inst_result_nxt[17]~19 (
	.dataa(!\A_ctrl_ld32~q ),
	.datab(!\d_readdata_d1[17]~q ),
	.datac(!\A_slow_ld_data_fill_bit~0_combout ),
	.datad(!src0_valid1),
	.datae(!q_a_17),
	.dataf(!\A_slow_inst_result_nxt[17]~30_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[17]~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[17]~19 .extended_lut = "off";
defparam \A_slow_inst_result_nxt[17]~19 .lut_mask = 64'h7FFFFFFFBFFFFFFF;
defparam \A_slow_inst_result_nxt[17]~19 .shared_arith = "off";

dffeas \A_slow_inst_result[17] (
	.clk(clk_clk),
	.d(\A_slow_inst_result_nxt[17]~19_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_ctrl_ld~q ),
	.q(\A_slow_inst_result[17]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[17] .is_wysiwyg = "true";
defparam \A_slow_inst_result[17] .power_up = "low";

cyclonev_lcell_comb \E_rot_mask[1]~1 (
	.dataa(!\E_src2[2]~q ),
	.datab(!\E_src2[1]~q ),
	.datac(!\E_src2[0]~q ),
	.datad(!\E_ctrl_shift_rot_right~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_mask[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_mask[1]~1 .extended_lut = "off";
defparam \E_rot_mask[1]~1 .lut_mask = 64'hFF7FFF7FFF7FFF7F;
defparam \E_rot_mask[1]~1 .shared_arith = "off";

dffeas \M_rot_mask[1] (
	.clk(clk_clk),
	.d(\E_rot_mask[1]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_rot_mask[1]~q ),
	.prn(vcc));
defparam \M_rot_mask[1] .is_wysiwyg = "true";
defparam \M_rot_mask[1] .power_up = "low";

cyclonev_lcell_comb \A_slow_inst_result_nxt[13]~45 (
	.dataa(!\d_readdata_d1[13]~q ),
	.datab(!\d_readdata_d1[29]~q ),
	.datac(!\A_slow_inst_result[9]~0_combout ),
	.datad(!\A_slow_inst_result[9]~1_combout ),
	.datae(!src0_valid),
	.dataf(!av_readdata_pre_13),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[13]~45_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[13]~45 .extended_lut = "off";
defparam \A_slow_inst_result_nxt[13]~45 .lut_mask = 64'h7FF7FFFFFFFFFFFF;
defparam \A_slow_inst_result_nxt[13]~45 .shared_arith = "off";

cyclonev_lcell_comb \A_slow_inst_result_nxt[13]~52 (
	.dataa(!\A_slow_inst_result_nxt[13]~45_combout ),
	.datab(!q_a_13),
	.datac(!\A_slow_ld_data_fill_bit~0_combout ),
	.datad(!src0_valid1),
	.datae(!\A_slow_inst_result[9]~0_combout ),
	.dataf(!\A_slow_inst_result[9]~1_combout ),
	.datag(!src_payload14),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[13]~52_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[13]~52 .extended_lut = "on";
defparam \A_slow_inst_result_nxt[13]~52 .lut_mask = 64'hFFD8FFD8FFD8FFD8;
defparam \A_slow_inst_result_nxt[13]~52 .shared_arith = "off";

dffeas \A_slow_inst_result[13] (
	.clk(clk_clk),
	.d(\A_slow_inst_result_nxt[13]~52_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_ctrl_ld~q ),
	.q(\A_slow_inst_result[13]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[13] .is_wysiwyg = "true";
defparam \A_slow_inst_result[13] .power_up = "low";

cyclonev_lcell_comb \A_slow_inst_result_nxt[9]~41 (
	.dataa(!\d_readdata_d1[9]~q ),
	.datab(!\d_readdata_d1[25]~q ),
	.datac(!\A_slow_inst_result[9]~0_combout ),
	.datad(!\A_slow_inst_result[9]~1_combout ),
	.datae(!src0_valid),
	.dataf(!av_readdata_pre_9),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[9]~41_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[9]~41 .extended_lut = "off";
defparam \A_slow_inst_result_nxt[9]~41 .lut_mask = 64'h7FF7FFFFFFFFFFFF;
defparam \A_slow_inst_result_nxt[9]~41 .shared_arith = "off";

cyclonev_lcell_comb \A_slow_inst_result_nxt[9]~64 (
	.dataa(!\A_slow_inst_result_nxt[9]~41_combout ),
	.datab(!q_a_9),
	.datac(!\A_slow_ld_data_fill_bit~0_combout ),
	.datad(!src0_valid1),
	.datae(!\A_slow_inst_result[9]~0_combout ),
	.dataf(!\A_slow_inst_result[9]~1_combout ),
	.datag(!src_payload8),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[9]~64_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[9]~64 .extended_lut = "on";
defparam \A_slow_inst_result_nxt[9]~64 .lut_mask = 64'hFFD8FFD8FFD8FFD8;
defparam \A_slow_inst_result_nxt[9]~64 .shared_arith = "off";

dffeas \A_slow_inst_result[9] (
	.clk(clk_clk),
	.d(\A_slow_inst_result_nxt[9]~64_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_ctrl_ld~q ),
	.q(\A_slow_inst_result[9]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[9] .is_wysiwyg = "true";
defparam \A_slow_inst_result[9] .power_up = "low";

dffeas \M_rot_prestep2[9] (
	.clk(clk_clk),
	.d(\E_rot_step1[5]~14_combout ),
	.asdata(\E_rot_step1[9]~15_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add10~1_combout ),
	.ena(!\A_mem_stall~q ),
	.q(\M_rot_prestep2[9]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[9] .is_wysiwyg = "true";
defparam \M_rot_prestep2[9] .power_up = "low";

cyclonev_lcell_comb \E_rot_step1[29]~8 (
	.dataa(!\E_src1[29]~q ),
	.datab(!\E_src1[28]~q ),
	.datac(!\E_src1[27]~q ),
	.datad(!\E_src1[26]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add10~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[29]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[29]~8 .extended_lut = "off";
defparam \E_rot_step1[29]~8 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[29]~8 .shared_arith = "off";

dffeas \M_rot_prestep2[1] (
	.clk(clk_clk),
	.d(\E_rot_step1[29]~8_combout ),
	.asdata(\E_rot_step1[1]~9_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add10~1_combout ),
	.ena(!\A_mem_stall~q ),
	.q(\M_rot_prestep2[1]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[1] .is_wysiwyg = "true";
defparam \M_rot_prestep2[1] .power_up = "low";

cyclonev_lcell_comb \A_slow_inst_result_nxt[19]~33 (
	.dataa(!\A_ctrl_ld32~q ),
	.datab(!\d_readdata_d1[19]~q ),
	.datac(!read_latency_shift_reg_01),
	.datad(!src0_valid),
	.datae(!av_readdata_pre_19),
	.dataf(!av_readdata_pre_191),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[19]~33_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[19]~33 .extended_lut = "off";
defparam \A_slow_inst_result_nxt[19]~33 .lut_mask = 64'h27FFFFFFFFFFFFFF;
defparam \A_slow_inst_result_nxt[19]~33 .shared_arith = "off";

cyclonev_lcell_comb \A_slow_inst_result_nxt[19]~18 (
	.dataa(!\A_ctrl_ld32~q ),
	.datab(!\A_ld_align_byte2_byte3_fill~q ),
	.datac(!\A_slow_ld_data_fill_bit~0_combout ),
	.datad(!src0_valid1),
	.datae(!q_a_19),
	.dataf(!\A_slow_inst_result_nxt[19]~33_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[19]~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[19]~18 .extended_lut = "off";
defparam \A_slow_inst_result_nxt[19]~18 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \A_slow_inst_result_nxt[19]~18 .shared_arith = "off";

dffeas \A_slow_inst_result[19] (
	.clk(clk_clk),
	.d(\A_slow_inst_result_nxt[19]~18_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_ctrl_ld~q ),
	.q(\A_slow_inst_result[19]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[19] .is_wysiwyg = "true";
defparam \A_slow_inst_result[19] .power_up = "low";

cyclonev_lcell_comb \E_rot_mask[3]~3 (
	.dataa(!\E_src2[2]~q ),
	.datab(!\E_src2[1]~q ),
	.datac(!\E_src2[0]~q ),
	.datad(!\E_ctrl_shift_rot_right~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_mask[3]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_mask[3]~3 .extended_lut = "off";
defparam \E_rot_mask[3]~3 .lut_mask = 64'hFF7FFF7FFF7FFF7F;
defparam \E_rot_mask[3]~3 .shared_arith = "off";

dffeas \M_rot_mask[3] (
	.clk(clk_clk),
	.d(\E_rot_mask[3]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_rot_mask[3]~q ),
	.prn(vcc));
defparam \M_rot_mask[3] .is_wysiwyg = "true";
defparam \M_rot_mask[3] .power_up = "low";

cyclonev_lcell_comb \A_slow_inst_result_nxt[15]~47 (
	.dataa(!\d_readdata_d1[15]~q ),
	.datab(!\d_readdata_d1[31]~q ),
	.datac(!\A_slow_inst_result[9]~0_combout ),
	.datad(!\A_slow_inst_result[9]~1_combout ),
	.datae(!src0_valid),
	.dataf(!av_readdata_pre_15),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[15]~47_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[15]~47 .extended_lut = "off";
defparam \A_slow_inst_result_nxt[15]~47 .lut_mask = 64'h7FF7FFFFFFFFFFFF;
defparam \A_slow_inst_result_nxt[15]~47 .shared_arith = "off";

cyclonev_lcell_comb \A_slow_inst_result_nxt[15]~60 (
	.dataa(!\A_slow_inst_result_nxt[15]~47_combout ),
	.datab(!q_a_15),
	.datac(!\A_slow_ld_data_fill_bit~0_combout ),
	.datad(!src0_valid1),
	.datae(!\A_slow_inst_result[9]~0_combout ),
	.dataf(!\A_slow_inst_result[9]~1_combout ),
	.datag(!src_payload12),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[15]~60_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[15]~60 .extended_lut = "on";
defparam \A_slow_inst_result_nxt[15]~60 .lut_mask = 64'hFFD8FFD8FFD8FFD8;
defparam \A_slow_inst_result_nxt[15]~60 .shared_arith = "off";

dffeas \A_slow_inst_result[15] (
	.clk(clk_clk),
	.d(\A_slow_inst_result_nxt[15]~60_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_ctrl_ld~q ),
	.q(\A_slow_inst_result[15]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[15] .is_wysiwyg = "true";
defparam \A_slow_inst_result[15] .power_up = "low";

cyclonev_lcell_comb \A_slow_inst_result_nxt[11]~43 (
	.dataa(!\d_readdata_d1[11]~q ),
	.datab(!\d_readdata_d1[27]~q ),
	.datac(!\A_slow_inst_result[9]~0_combout ),
	.datad(!\A_slow_inst_result[9]~1_combout ),
	.datae(!src0_valid),
	.dataf(!av_readdata_pre_11),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[11]~43_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[11]~43 .extended_lut = "off";
defparam \A_slow_inst_result_nxt[11]~43 .lut_mask = 64'h7FF7FFFFFFFFFFFF;
defparam \A_slow_inst_result_nxt[11]~43 .shared_arith = "off";

cyclonev_lcell_comb \A_slow_inst_result_nxt[11]~76 (
	.dataa(!\A_slow_inst_result[9]~1_combout ),
	.datab(!\A_slow_inst_result_nxt[11]~43_combout ),
	.datac(!\A_slow_ld_data_fill_bit~0_combout ),
	.datad(!src_payload5),
	.datae(!\A_slow_inst_result[9]~0_combout ),
	.dataf(!q_a_11),
	.datag(!src0_valid1),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[11]~76_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[11]~76 .extended_lut = "on";
defparam \A_slow_inst_result_nxt[11]~76 .lut_mask = 64'hFFD8FFD8FFD8FFD8;
defparam \A_slow_inst_result_nxt[11]~76 .shared_arith = "off";

dffeas \A_slow_inst_result[11] (
	.clk(clk_clk),
	.d(\A_slow_inst_result_nxt[11]~76_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_ctrl_ld~q ),
	.q(\A_slow_inst_result[11]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[11] .is_wysiwyg = "true";
defparam \A_slow_inst_result[11] .power_up = "low";

dffeas \M_rot_prestep2[11] (
	.clk(clk_clk),
	.d(\E_rot_step1[7]~30_combout ),
	.asdata(\E_rot_step1[11]~31_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add10~1_combout ),
	.ena(!\A_mem_stall~q ),
	.q(\M_rot_prestep2[11]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[11] .is_wysiwyg = "true";
defparam \M_rot_prestep2[11] .power_up = "low";

cyclonev_lcell_comb \E_rot_step1[31]~24 (
	.dataa(!\E_src1[31]~q ),
	.datab(!\E_src1[30]~q ),
	.datac(!\E_src1[29]~q ),
	.datad(!\E_src1[28]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add10~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[31]~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[31]~24 .extended_lut = "off";
defparam \E_rot_step1[31]~24 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[31]~24 .shared_arith = "off";

dffeas \M_rot_prestep2[3] (
	.clk(clk_clk),
	.d(\E_rot_step1[31]~24_combout ),
	.asdata(\E_rot_step1[3]~25_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add10~1_combout ),
	.ena(!\A_mem_stall~q ),
	.q(\M_rot_prestep2[3]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[3] .is_wysiwyg = "true";
defparam \M_rot_prestep2[3] .power_up = "low";

cyclonev_lcell_comb \E_rot_step1[23]~26 (
	.dataa(!\E_src1[23]~q ),
	.datab(!\E_src1[22]~q ),
	.datac(!\E_src1[21]~q ),
	.datad(!\E_src1[20]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add10~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[23]~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[23]~26 .extended_lut = "off";
defparam \E_rot_step1[23]~26 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[23]~26 .shared_arith = "off";

cyclonev_lcell_comb \E_rot_step1[27]~27 (
	.dataa(!\E_src1[27]~q ),
	.datab(!\E_src1[26]~q ),
	.datac(!\E_src1[25]~q ),
	.datad(!\E_src1[24]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add10~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[27]~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[27]~27 .extended_lut = "off";
defparam \E_rot_step1[27]~27 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[27]~27 .shared_arith = "off";

dffeas \M_rot_prestep2[27] (
	.clk(clk_clk),
	.d(\E_rot_step1[23]~26_combout ),
	.asdata(\E_rot_step1[27]~27_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add10~1_combout ),
	.ena(!\A_mem_stall~q ),
	.q(\M_rot_prestep2[27]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[27] .is_wysiwyg = "true";
defparam \M_rot_prestep2[27] .power_up = "low";

cyclonev_lcell_comb \Add10~2 (
	.dataa(!\E_src2[3]~q ),
	.datab(!\E_src2[2]~q ),
	.datac(!\E_src2[1]~q ),
	.datad(!\E_src2[0]~q ),
	.datae(!\E_ctrl_shift_rot_right~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add10~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add10~2 .extended_lut = "off";
defparam \Add10~2 .lut_mask = 64'h9669699696696996;
defparam \Add10~2 .shared_arith = "off";

dffeas \M_rot_rn[3] (
	.clk(clk_clk),
	.d(\Add10~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_rot_rn[3]~q ),
	.prn(vcc));
defparam \M_rot_rn[3] .is_wysiwyg = "true";
defparam \M_rot_rn[3] .power_up = "low";

cyclonev_lcell_comb \Add10~3 (
	.dataa(!\E_src2[3]~q ),
	.datab(!\E_src2[2]~q ),
	.datac(!\E_src2[1]~q ),
	.datad(!\E_src2[0]~q ),
	.datae(!\E_src2[4]~q ),
	.dataf(!\E_ctrl_shift_rot_right~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add10~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add10~3 .extended_lut = "off";
defparam \Add10~3 .lut_mask = 64'h6996966996696996;
defparam \Add10~3 .shared_arith = "off";

dffeas \M_rot_rn[4] (
	.clk(clk_clk),
	.d(\Add10~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_rot_rn[4]~q ),
	.prn(vcc));
defparam \M_rot_rn[4] .is_wysiwyg = "true";
defparam \M_rot_rn[4] .power_up = "low";

cyclonev_lcell_comb \M_rot[3]~14 (
	.dataa(!\M_rot_prestep2[11]~q ),
	.datab(!\M_rot_prestep2[3]~q ),
	.datac(!\M_rot_prestep2[27]~q ),
	.datad(!\M_rot_prestep2[19]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[3]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[3]~14 .extended_lut = "off";
defparam \M_rot[3]~14 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[3]~14 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~14 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_mask[3]~q ),
	.datac(!\M_rot_pass1~q ),
	.datad(!\M_rot_sel_fill1~q ),
	.datae(!\M_rot[3]~14_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~14 .extended_lut = "off";
defparam \A_shift_rot_result~14 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~14 .shared_arith = "off";

dffeas \A_shift_rot_result[11] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~14_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_shift_rot_result[11]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[11] .is_wysiwyg = "true";
defparam \A_shift_rot_result[11] .power_up = "low";

dffeas \E_pc[9] (
	.clk(clk_clk),
	.d(\D_pc[9]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_pc[9]~q ),
	.prn(vcc));
defparam \E_pc[9] .is_wysiwyg = "true";
defparam \E_pc[9] .power_up = "low";

dffeas \E_pc[8] (
	.clk(clk_clk),
	.d(\D_pc[8]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_pc[8]~q ),
	.prn(vcc));
defparam \E_pc[8] .is_wysiwyg = "true";
defparam \E_pc[8] .power_up = "low";

dffeas \E_pc[7] (
	.clk(clk_clk),
	.d(\D_pc[7]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_pc[7]~q ),
	.prn(vcc));
defparam \E_pc[7] .is_wysiwyg = "true";
defparam \E_pc[7] .power_up = "low";

dffeas \E_pc[6] (
	.clk(clk_clk),
	.d(\D_pc[6]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_pc[6]~q ),
	.prn(vcc));
defparam \E_pc[6] .is_wysiwyg = "true";
defparam \E_pc[6] .power_up = "low";

cyclonev_lcell_comb \Add7~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_pc[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add7~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add7~29_sumout ),
	.cout(\Add7~30 ),
	.shareout());
defparam \Add7~29 .extended_lut = "off";
defparam \Add7~29 .lut_mask = 64'h00000000000000FF;
defparam \Add7~29 .shared_arith = "off";

cyclonev_lcell_comb \Add7~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_pc[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add7~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add7~33_sumout ),
	.cout(\Add7~34 ),
	.shareout());
defparam \Add7~33 .extended_lut = "off";
defparam \Add7~33 .lut_mask = 64'h00000000000000FF;
defparam \Add7~33 .shared_arith = "off";

cyclonev_lcell_comb \Add7~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_pc[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add7~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add7~25_sumout ),
	.cout(\Add7~26 ),
	.shareout());
defparam \Add7~25 .extended_lut = "off";
defparam \Add7~25 .lut_mask = 64'h00000000000000FF;
defparam \Add7~25 .shared_arith = "off";

cyclonev_lcell_comb \Add7~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_pc[9]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add7~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add7~21_sumout ),
	.cout(\Add7~22 ),
	.shareout());
defparam \Add7~21 .extended_lut = "off";
defparam \Add7~21 .lut_mask = 64'h00000000000000FF;
defparam \Add7~21 .shared_arith = "off";

dffeas \M_pc_plus_one[9] (
	.clk(clk_clk),
	.d(\Add7~21_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_pc_plus_one[9]~q ),
	.prn(vcc));
defparam \M_pc_plus_one[9] .is_wysiwyg = "true";
defparam \M_pc_plus_one[9] .power_up = "low";

cyclonev_lcell_comb \E_op_rdctl~1 (
	.dataa(!\E_iw[15]~q ),
	.datab(!\E_iw[12]~q ),
	.datac(!\E_op_rdctl~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_op_rdctl~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_op_rdctl~1 .extended_lut = "off";
defparam \E_op_rdctl~1 .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \E_op_rdctl~1 .shared_arith = "off";

cyclonev_lcell_comb E_op_rdctl(
	.dataa(!\E_iw[14]~q ),
	.datab(!\E_op_rdctl~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_op_rdctl~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam E_op_rdctl.extended_lut = "off";
defparam E_op_rdctl.lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam E_op_rdctl.shared_arith = "off";

dffeas M_ctrl_rd_ctl_reg(
	.clk(clk_clk),
	.d(\E_op_rdctl~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_ctrl_rd_ctl_reg~q ),
	.prn(vcc));
defparam M_ctrl_rd_ctl_reg.is_wysiwyg = "true";
defparam M_ctrl_rd_ctl_reg.power_up = "low";

cyclonev_lcell_comb \A_inst_result[9]~0 (
	.dataa(!\M_exc_any~combout ),
	.datab(!\M_ctrl_rd_ctl_reg~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_inst_result[9]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_inst_result[9]~0 .extended_lut = "off";
defparam \A_inst_result[9]~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \A_inst_result[9]~0 .shared_arith = "off";

dffeas \A_inst_result[11] (
	.clk(clk_clk),
	.d(\M_pc_plus_one[9]~q ),
	.asdata(\M_alu_result[11]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\A_inst_result[9]~0_combout ),
	.sload(!\M_exc_any~combout ),
	.ena(!\A_mem_stall~q ),
	.q(\A_inst_result[11]~q ),
	.prn(vcc));
defparam \A_inst_result[11] .is_wysiwyg = "true";
defparam \A_inst_result[11] .power_up = "low";

dffeas \A_mul_cell_p1[11] (
	.clk(clk_clk),
	.d(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[11]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_mul_cell_p1[11]~q ),
	.prn(vcc));
defparam \A_mul_cell_p1[11] .is_wysiwyg = "true";
defparam \A_mul_cell_p1[11] .power_up = "low";

cyclonev_lcell_comb \Equal95~7 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[1]~q ),
	.datac(!\D_iw[2]~q ),
	.datad(!\D_iw[3]~q ),
	.datae(!\D_iw[4]~q ),
	.dataf(!\D_iw[5]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal95~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal95~7 .extended_lut = "off";
defparam \Equal95~7 .lut_mask = 64'hFFFFFFEFFFFFFFFF;
defparam \Equal95~7 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_late_result~2 (
	.dataa(!\D_iw[16]~q ),
	.datab(!\D_iw[13]~q ),
	.datac(!\D_iw[12]~q ),
	.datad(!\D_iw[11]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_late_result~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_late_result~2 .extended_lut = "off";
defparam \D_ctrl_late_result~2 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \D_ctrl_late_result~2 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_mul_lsw~0 (
	.dataa(!\Equal95~0_combout ),
	.datab(!\Equal95~7_combout ),
	.datac(!\D_ctrl_late_result~2_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_mul_lsw~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_mul_lsw~0 .extended_lut = "off";
defparam \D_ctrl_mul_lsw~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \D_ctrl_mul_lsw~0 .shared_arith = "off";

dffeas E_ctrl_mul_lsw(
	.clk(clk_clk),
	.d(\D_ctrl_mul_lsw~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_ctrl_mul_lsw~q ),
	.prn(vcc));
defparam E_ctrl_mul_lsw.is_wysiwyg = "true";
defparam E_ctrl_mul_lsw.power_up = "low";

dffeas M_ctrl_mul_lsw(
	.clk(clk_clk),
	.d(\E_ctrl_mul_lsw~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_ctrl_mul_lsw~q ),
	.prn(vcc));
defparam M_ctrl_mul_lsw.is_wysiwyg = "true";
defparam M_ctrl_mul_lsw.power_up = "low";

dffeas A_ctrl_mul_lsw(
	.clk(clk_clk),
	.d(\M_ctrl_mul_lsw~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_ctrl_mul_lsw~q ),
	.prn(vcc));
defparam A_ctrl_mul_lsw.is_wysiwyg = "true";
defparam A_ctrl_mul_lsw.power_up = "low";

cyclonev_lcell_comb \D_ctrl_shift_rot~0 (
	.dataa(!\Equal95~0_combout ),
	.datab(!\D_iw[13]~q ),
	.datac(!\D_iw[12]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_shift_rot~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_shift_rot~0 .extended_lut = "off";
defparam \D_ctrl_shift_rot~0 .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \D_ctrl_shift_rot~0 .shared_arith = "off";

dffeas E_ctrl_shift_rot(
	.clk(clk_clk),
	.d(\D_ctrl_shift_rot~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_ctrl_shift_rot~q ),
	.prn(vcc));
defparam E_ctrl_shift_rot.is_wysiwyg = "true";
defparam E_ctrl_shift_rot.power_up = "low";

dffeas M_ctrl_shift_rot(
	.clk(clk_clk),
	.d(\E_ctrl_shift_rot~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_ctrl_shift_rot~q ),
	.prn(vcc));
defparam M_ctrl_shift_rot.is_wysiwyg = "true";
defparam M_ctrl_shift_rot.power_up = "low";

dffeas A_ctrl_shift_rot(
	.clk(clk_clk),
	.d(\M_ctrl_shift_rot~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_ctrl_shift_rot~q ),
	.prn(vcc));
defparam A_ctrl_shift_rot.is_wysiwyg = "true";
defparam A_ctrl_shift_rot.power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[15]~0 (
	.dataa(!\A_exc_any~q ),
	.datab(!\A_ctrl_mul_lsw~q ),
	.datac(!\A_ctrl_shift_rot~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[15]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[15]~0 .extended_lut = "off";
defparam \A_wr_data_unfiltered[15]~0 .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \A_wr_data_unfiltered[15]~0 .shared_arith = "off";

cyclonev_lcell_comb \A_slow_inst_sel_nxt~0 (
	.dataa(!\A_mem_stall~q ),
	.datab(!\A_ctrl_ld~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_sel_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_sel_nxt~0 .extended_lut = "off";
defparam \A_slow_inst_sel_nxt~0 .lut_mask = 64'h7777777777777777;
defparam \A_slow_inst_sel_nxt~0 .shared_arith = "off";

dffeas A_slow_inst_sel(
	.clk(clk_clk),
	.d(\A_slow_inst_sel_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_slow_inst_sel~q ),
	.prn(vcc));
defparam A_slow_inst_sel.is_wysiwyg = "true";
defparam A_slow_inst_sel.power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[15]~1 (
	.dataa(!\A_exc_any~q ),
	.datab(!\A_ctrl_mul_lsw~q ),
	.datac(!\A_ctrl_shift_rot~q ),
	.datad(!\A_slow_inst_sel~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[15]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[15]~1 .extended_lut = "off";
defparam \A_wr_data_unfiltered[15]~1 .lut_mask = 64'hEFFFEFFFEFFFEFFF;
defparam \A_wr_data_unfiltered[15]~1 .shared_arith = "off";

cyclonev_lcell_comb \A_wr_data_unfiltered[11]~16 (
	.dataa(!\A_slow_inst_result[11]~q ),
	.datab(!\A_shift_rot_result[11]~q ),
	.datac(!\A_inst_result[11]~q ),
	.datad(!\A_mul_cell_p1[11]~q ),
	.datae(!\A_wr_data_unfiltered[15]~0_combout ),
	.dataf(!\A_wr_data_unfiltered[15]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[11]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[11]~16 .extended_lut = "off";
defparam \A_wr_data_unfiltered[11]~16 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_wr_data_unfiltered[11]~16 .shared_arith = "off";

dffeas \W_wr_data[11] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[11]~16_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[11]~q ),
	.prn(vcc));
defparam \W_wr_data[11] .is_wysiwyg = "true";
defparam \W_wr_data[11] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[11]~38 (
	.dataa(!\D_src2_reg[0]~7_combout ),
	.datab(!\D_src2_reg[0]~8_combout ),
	.datac(!\W_wr_data[11]~q ),
	.datad(!\A_wr_data_unfiltered[11]~16_combout ),
	.datae(!\M_alu_result[11]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[11]~38_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[11]~38 .extended_lut = "off";
defparam \D_src2_reg[11]~38 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \D_src2_reg[11]~38 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[11]~39 (
	.dataa(!\D_src2_reg[0]~4_combout ),
	.datab(!\D_src2_reg[0]~5_combout ),
	.datac(!\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[11] ),
	.datad(!\E_alu_result[11]~combout ),
	.datae(!\D_src2_reg[11]~38_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[11]~39_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[11]~39 .extended_lut = "off";
defparam \D_src2_reg[11]~39 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \D_src2_reg[11]~39 .shared_arith = "off";

cyclonev_lcell_comb \E_src2[5]~2 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\D_ctrl_src2_choose_imm~q ),
	.datac(!\D_ctrl_hi_imm16~q ),
	.datad(!\D_ctrl_shift_right_arith~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_src2[5]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_src2[5]~2 .extended_lut = "off";
defparam \E_src2[5]~2 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \E_src2[5]~2 .shared_arith = "off";

dffeas \E_src2[11] (
	.clk(clk_clk),
	.d(\D_iw[17]~q ),
	.asdata(\D_src2_reg[11]~39_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src2[5]~2_combout ),
	.sload(!\D_ctrl_src2_choose_imm~q ),
	.ena(!\A_mem_stall~q ),
	.q(\E_src2[11]~q ),
	.prn(vcc));
defparam \E_src2[11] .is_wysiwyg = "true";
defparam \E_src2[11] .power_up = "low";

cyclonev_lcell_comb \Add9~45 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[7]~q ),
	.datae(gnd),
	.dataf(!\E_src1[7]~q ),
	.datag(gnd),
	.cin(\Add9~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~45_sumout ),
	.cout(\Add9~46 ),
	.shareout());
defparam \Add9~45 .extended_lut = "off";
defparam \Add9~45 .lut_mask = 64'h0000FF00000055AA;
defparam \Add9~45 .shared_arith = "off";

cyclonev_lcell_comb \Add9~9 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[8]~q ),
	.datae(gnd),
	.dataf(!\E_src1[8]~q ),
	.datag(gnd),
	.cin(\Add9~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~9_sumout ),
	.cout(\Add9~10 ),
	.shareout());
defparam \Add9~9 .extended_lut = "off";
defparam \Add9~9 .lut_mask = 64'h0000FF00000055AA;
defparam \Add9~9 .shared_arith = "off";

cyclonev_lcell_comb \Add9~41 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[9]~q ),
	.datae(gnd),
	.dataf(!\E_src1[9]~q ),
	.datag(gnd),
	.cin(\Add9~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~41_sumout ),
	.cout(\Add9~42 ),
	.shareout());
defparam \Add9~41 .extended_lut = "off";
defparam \Add9~41 .lut_mask = 64'h0000FF00000055AA;
defparam \Add9~41 .shared_arith = "off";

cyclonev_lcell_comb \Add9~37 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[10]~q ),
	.datae(gnd),
	.dataf(!\E_src1[10]~q ),
	.datag(gnd),
	.cin(\Add9~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~37_sumout ),
	.cout(\Add9~38 ),
	.shareout());
defparam \Add9~37 .extended_lut = "off";
defparam \Add9~37 .lut_mask = 64'h0000FF00000055AA;
defparam \Add9~37 .shared_arith = "off";

cyclonev_lcell_comb \Add9~33 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[11]~q ),
	.datae(gnd),
	.dataf(!\E_src1[11]~q ),
	.datag(gnd),
	.cin(\Add9~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~33_sumout ),
	.cout(\Add9~34 ),
	.shareout());
defparam \Add9~33 .extended_lut = "off";
defparam \Add9~33 .lut_mask = 64'h0000FF00000055AA;
defparam \Add9~33 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result~11 (
	.dataa(!\E_src2[11]~q ),
	.datab(!\E_src1[11]~q ),
	.datac(!\E_logic_op[1]~q ),
	.datad(!\E_logic_op[0]~q ),
	.datae(!\E_ctrl_logic~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result~11 .extended_lut = "off";
defparam \E_alu_result~11 .lut_mask = 64'h6996FFFF6996FFFF;
defparam \E_alu_result~11 .shared_arith = "off";

dffeas \D_pc_plus_one[9] (
	.clk(clk_clk),
	.d(\Add3~41_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_pc_plus_one[9]~q ),
	.prn(vcc));
defparam \D_pc_plus_one[9] .is_wysiwyg = "true";
defparam \D_pc_plus_one[9] .power_up = "low";

dffeas \E_extra_pc[9] (
	.clk(clk_clk),
	.d(\D_br_taken_waddr_partial[9]~q ),
	.asdata(\D_pc_plus_one[9]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_br_pred_not_taken~combout ),
	.ena(!\A_mem_stall~q ),
	.q(\E_extra_pc[9]~q ),
	.prn(vcc));
defparam \E_extra_pc[9] .is_wysiwyg = "true";
defparam \E_extra_pc[9] .power_up = "low";

cyclonev_lcell_comb \E_alu_result[11] (
	.dataa(!\Add9~33_sumout ),
	.datab(!\E_ctrl_retaddr~q ),
	.datac(!\E_alu_result~0_combout ),
	.datad(!\E_alu_result~11_combout ),
	.datae(!\E_extra_pc[9]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[11]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[11] .extended_lut = "off";
defparam \E_alu_result[11] .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \E_alu_result[11] .shared_arith = "off";

dffeas \M_alu_result[11] (
	.clk(clk_clk),
	.d(\E_alu_result[11]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_alu_result[11]~q ),
	.prn(vcc));
defparam \M_alu_result[11] .is_wysiwyg = "true";
defparam \M_alu_result[11] .power_up = "low";

cyclonev_lcell_comb \F_ctrl_a_not_src~0 (
	.dataa(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[1] ),
	.datab(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[2] ),
	.datac(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[3] ),
	.datad(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[4] ),
	.datae(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[5] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ctrl_a_not_src~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ctrl_a_not_src~0 .extended_lut = "off";
defparam \F_ctrl_a_not_src~0 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \F_ctrl_a_not_src~0 .shared_arith = "off";

dffeas D_ctrl_a_not_src(
	.clk(clk_clk),
	.d(\F_ctrl_a_not_src~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_ctrl_a_not_src~q ),
	.prn(vcc));
defparam D_ctrl_a_not_src.is_wysiwyg = "true";
defparam D_ctrl_a_not_src.power_up = "low";

cyclonev_lcell_comb \E_regnum_a_cmp_F~0 (
	.dataa(!\E_wr_dst_reg~combout ),
	.datab(!\E_dst_regnum[0]~q ),
	.datac(!\E_dst_regnum[1]~q ),
	.datad(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[27] ),
	.datae(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[28] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_regnum_a_cmp_F~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_regnum_a_cmp_F~0 .extended_lut = "off";
defparam \E_regnum_a_cmp_F~0 .lut_mask = 64'h7DD7D77D7DD7D77D;
defparam \E_regnum_a_cmp_F~0 .shared_arith = "off";

cyclonev_lcell_comb \E_regnum_a_cmp_F~1 (
	.dataa(!\E_dst_regnum[2]~q ),
	.datab(!\E_dst_regnum[3]~q ),
	.datac(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[29] ),
	.datad(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[30] ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_regnum_a_cmp_F~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_regnum_a_cmp_F~1 .extended_lut = "off";
defparam \E_regnum_a_cmp_F~1 .lut_mask = 64'h6996699669966996;
defparam \E_regnum_a_cmp_F~1 .shared_arith = "off";

cyclonev_lcell_comb E_regnum_a_cmp_F(
	.dataa(!\E_dst_regnum[4]~q ),
	.datab(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[31] ),
	.datac(!\E_regnum_a_cmp_F~0_combout ),
	.datad(!\E_regnum_a_cmp_F~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_regnum_a_cmp_F~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam E_regnum_a_cmp_F.extended_lut = "off";
defparam E_regnum_a_cmp_F.lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam E_regnum_a_cmp_F.shared_arith = "off";

cyclonev_lcell_comb \D_regnum_a_cmp_F~0 (
	.dataa(!\D_dst_regnum[0]~2_combout ),
	.datab(!\D_dst_regnum[2]~3_combout ),
	.datac(!\D_dst_regnum[3]~4_combout ),
	.datad(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[27] ),
	.datae(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[29] ),
	.dataf(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[30] ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_regnum_a_cmp_F~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_regnum_a_cmp_F~0 .extended_lut = "off";
defparam \D_regnum_a_cmp_F~0 .lut_mask = 64'h6996966996696996;
defparam \D_regnum_a_cmp_F~0 .shared_arith = "off";

cyclonev_lcell_comb D_regnum_a_cmp_F(
	.dataa(!\D_dst_regnum[1]~0_combout ),
	.datab(!\D_dst_regnum[4]~1_combout ),
	.datac(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[28] ),
	.datad(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[31] ),
	.datae(!\D_wr_dst_reg~combout ),
	.dataf(!\D_regnum_a_cmp_F~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_regnum_a_cmp_F~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam D_regnum_a_cmp_F.extended_lut = "off";
defparam D_regnum_a_cmp_F.lut_mask = 64'h6996FFFFFFFFFFFF;
defparam D_regnum_a_cmp_F.shared_arith = "off";

dffeas E_regnum_a_cmp_D(
	.clk(clk_clk),
	.d(\D_regnum_a_cmp_F~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\F_stall~0_combout ),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_regnum_a_cmp_D~q ),
	.prn(vcc));
defparam E_regnum_a_cmp_D.is_wysiwyg = "true";
defparam E_regnum_a_cmp_D.power_up = "low";

dffeas M_regnum_a_cmp_D(
	.clk(clk_clk),
	.d(\E_regnum_a_cmp_F~combout ),
	.asdata(\E_regnum_a_cmp_D~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\F_stall~0_combout ),
	.ena(!\A_mem_stall~q ),
	.q(\M_regnum_a_cmp_D~q ),
	.prn(vcc));
defparam M_regnum_a_cmp_D.is_wysiwyg = "true";
defparam M_regnum_a_cmp_D.power_up = "low";

cyclonev_lcell_comb \A_regnum_a_cmp_F~0 (
	.dataa(!\A_dst_regnum~1_combout ),
	.datab(!\A_dst_regnum~2_combout ),
	.datac(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[28] ),
	.datad(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[29] ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_regnum_a_cmp_F~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_regnum_a_cmp_F~0 .extended_lut = "off";
defparam \A_regnum_a_cmp_F~0 .lut_mask = 64'h6996699669966996;
defparam \A_regnum_a_cmp_F~0 .shared_arith = "off";

cyclonev_lcell_comb \A_regnum_a_cmp_F~1 (
	.dataa(!\A_dst_regnum~3_combout ),
	.datab(!\A_dst_regnum~4_combout ),
	.datac(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[30] ),
	.datad(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[31] ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_regnum_a_cmp_F~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_regnum_a_cmp_F~1 .extended_lut = "off";
defparam \A_regnum_a_cmp_F~1 .lut_mask = 64'h6996699669966996;
defparam \A_regnum_a_cmp_F~1 .shared_arith = "off";

cyclonev_lcell_comb A_regnum_a_cmp_F(
	.dataa(!\A_wr_dst_reg~0_combout ),
	.datab(!\A_dst_regnum~0_combout ),
	.datac(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[27] ),
	.datad(!\A_regnum_a_cmp_F~0_combout ),
	.datae(!\A_regnum_a_cmp_F~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_regnum_a_cmp_F~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam A_regnum_a_cmp_F.extended_lut = "off";
defparam A_regnum_a_cmp_F.lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam A_regnum_a_cmp_F.shared_arith = "off";

cyclonev_lcell_comb \M_regnum_a_cmp_F~0 (
	.dataa(!\M_dst_regnum[0]~q ),
	.datab(!\M_dst_regnum[1]~q ),
	.datac(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[27] ),
	.datad(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[28] ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_regnum_a_cmp_F~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_regnum_a_cmp_F~0 .extended_lut = "off";
defparam \M_regnum_a_cmp_F~0 .lut_mask = 64'h6996699669966996;
defparam \M_regnum_a_cmp_F~0 .shared_arith = "off";

cyclonev_lcell_comb \M_regnum_a_cmp_F~1 (
	.dataa(!\M_dst_regnum[3]~q ),
	.datab(!\M_dst_regnum[4]~q ),
	.datac(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[30] ),
	.datad(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[31] ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_regnum_a_cmp_F~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_regnum_a_cmp_F~1 .extended_lut = "off";
defparam \M_regnum_a_cmp_F~1 .lut_mask = 64'h6996699669966996;
defparam \M_regnum_a_cmp_F~1 .shared_arith = "off";

cyclonev_lcell_comb M_regnum_a_cmp_F(
	.dataa(!\M_dst_regnum[2]~q ),
	.datab(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[29] ),
	.datac(!\M_wr_dst_reg~0_combout ),
	.datad(!\M_regnum_a_cmp_F~0_combout ),
	.datae(!\M_regnum_a_cmp_F~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_regnum_a_cmp_F~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam M_regnum_a_cmp_F.extended_lut = "off";
defparam M_regnum_a_cmp_F.lut_mask = 64'hF6FFFFFFF6FFFFFF;
defparam M_regnum_a_cmp_F.shared_arith = "off";

dffeas A_regnum_a_cmp_D(
	.clk(clk_clk),
	.d(\M_regnum_a_cmp_F~combout ),
	.asdata(\M_regnum_a_cmp_D~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\F_stall~0_combout ),
	.ena(!\A_mem_stall~q ),
	.q(\A_regnum_a_cmp_D~q ),
	.prn(vcc));
defparam A_regnum_a_cmp_D.is_wysiwyg = "true";
defparam A_regnum_a_cmp_D.power_up = "low";

dffeas W_regnum_a_cmp_D(
	.clk(clk_clk),
	.d(\A_regnum_a_cmp_F~combout ),
	.asdata(\A_regnum_a_cmp_D~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\F_stall~0_combout ),
	.ena(vcc),
	.q(\W_regnum_a_cmp_D~q ),
	.prn(vcc));
defparam W_regnum_a_cmp_D.is_wysiwyg = "true";
defparam W_regnum_a_cmp_D.power_up = "low";

cyclonev_lcell_comb \E_src1[26]~0 (
	.dataa(!\D_ctrl_a_not_src~q ),
	.datab(!\M_regnum_a_cmp_D~q ),
	.datac(!\W_regnum_a_cmp_D~q ),
	.datad(!\A_regnum_a_cmp_D~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_src1[26]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_src1[26]~0 .extended_lut = "off";
defparam \E_src1[26]~0 .lut_mask = 64'hEFFFEFFFEFFFEFFF;
defparam \E_src1[26]~0 .shared_arith = "off";

cyclonev_lcell_comb \E_src1[26]~1 (
	.dataa(!\D_ctrl_a_not_src~q ),
	.datab(!\M_regnum_a_cmp_D~q ),
	.datac(!\A_regnum_a_cmp_D~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_src1[26]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_src1[26]~1 .extended_lut = "off";
defparam \E_src1[26]~1 .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \E_src1[26]~1 .shared_arith = "off";

cyclonev_lcell_comb \D_src1_reg[11]~10 (
	.dataa(!\M_alu_result[11]~q ),
	.datab(!\A_wr_data_unfiltered[11]~16_combout ),
	.datac(!\first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[11] ),
	.datad(!\W_wr_data[11]~q ),
	.datae(!\E_src1[26]~0_combout ),
	.dataf(!\E_src1[26]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[11]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[11]~10 .extended_lut = "off";
defparam \D_src1_reg[11]~10 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[11]~10 .shared_arith = "off";

dffeas \D_iw[31] (
	.clk(clk_clk),
	.d(\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[31] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_iw[31]~q ),
	.prn(vcc));
defparam \D_iw[31] .is_wysiwyg = "true";
defparam \D_iw[31] .power_up = "low";

dffeas \D_iw[30] (
	.clk(clk_clk),
	.d(\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[30] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_iw[30]~q ),
	.prn(vcc));
defparam \D_iw[30] .is_wysiwyg = "true";
defparam \D_iw[30] .power_up = "low";

dffeas \D_iw[29] (
	.clk(clk_clk),
	.d(\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[29] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_iw[29]~q ),
	.prn(vcc));
defparam \D_iw[29] .is_wysiwyg = "true";
defparam \D_iw[29] .power_up = "low";

dffeas \D_iw[28] (
	.clk(clk_clk),
	.d(\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[28] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_iw[28]~q ),
	.prn(vcc));
defparam \D_iw[28] .is_wysiwyg = "true";
defparam \D_iw[28] .power_up = "low";

dffeas \D_iw[27] (
	.clk(clk_clk),
	.d(\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[27] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_iw[27]~q ),
	.prn(vcc));
defparam \D_iw[27] .is_wysiwyg = "true";
defparam \D_iw[27] .power_up = "low";

cyclonev_lcell_comb \Equal303~0 (
	.dataa(!\D_iw[31]~q ),
	.datab(!\D_iw[30]~q ),
	.datac(!\D_iw[29]~q ),
	.datad(!\D_iw[28]~q ),
	.datae(!\D_iw[27]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal303~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal303~0 .extended_lut = "off";
defparam \Equal303~0 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \Equal303~0 .shared_arith = "off";

cyclonev_lcell_comb D_src1_hazard_E(
	.dataa(!\D_ctrl_a_not_src~q ),
	.datab(!\E_regnum_a_cmp_D~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_hazard_E~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam D_src1_hazard_E.extended_lut = "off";
defparam D_src1_hazard_E.lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam D_src1_hazard_E.shared_arith = "off";

dffeas \E_src1[11] (
	.clk(clk_clk),
	.d(\D_src1_reg[11]~10_combout ),
	.asdata(\E_alu_result[11]~combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\Equal303~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(!\A_mem_stall~q ),
	.q(\E_src1[11]~q ),
	.prn(vcc));
defparam \E_src1[11] .is_wysiwyg = "true";
defparam \E_src1[11] .power_up = "low";

cyclonev_lcell_comb \E_rot_step1[11]~31 (
	.dataa(!\E_src1[11]~q ),
	.datab(!\E_src1[10]~q ),
	.datac(!\E_src1[9]~q ),
	.datad(!\E_src1[8]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add10~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[11]~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[11]~31 .extended_lut = "off";
defparam \E_rot_step1[11]~31 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[11]~31 .shared_arith = "off";

dffeas \M_rot_prestep2[15] (
	.clk(clk_clk),
	.d(\E_rot_step1[11]~31_combout ),
	.asdata(\E_rot_step1[15]~28_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add10~1_combout ),
	.ena(!\A_mem_stall~q ),
	.q(\M_rot_prestep2[15]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[15] .is_wysiwyg = "true";
defparam \M_rot_prestep2[15] .power_up = "low";

dffeas \M_rot_prestep2[31] (
	.clk(clk_clk),
	.d(\E_rot_step1[27]~27_combout ),
	.asdata(\E_rot_step1[31]~24_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add10~1_combout ),
	.ena(!\A_mem_stall~q ),
	.q(\M_rot_prestep2[31]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[31] .is_wysiwyg = "true";
defparam \M_rot_prestep2[31] .power_up = "low";

cyclonev_lcell_comb \E_rot_step1[19]~29 (
	.dataa(!\E_src1[19]~q ),
	.datab(!\E_src1[18]~q ),
	.datac(!\E_src1[17]~q ),
	.datad(!\E_src1[16]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add10~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[19]~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[19]~29 .extended_lut = "off";
defparam \E_rot_step1[19]~29 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[19]~29 .shared_arith = "off";

dffeas \M_rot_prestep2[23] (
	.clk(clk_clk),
	.d(\E_rot_step1[19]~29_combout ),
	.asdata(\E_rot_step1[23]~26_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add10~1_combout ),
	.ena(!\A_mem_stall~q ),
	.q(\M_rot_prestep2[23]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[23] .is_wysiwyg = "true";
defparam \M_rot_prestep2[23] .power_up = "low";

cyclonev_lcell_comb \M_rot[7]~27 (
	.dataa(!\M_rot_prestep2[15]~q ),
	.datab(!\M_rot_prestep2[7]~q ),
	.datac(!\M_rot_prestep2[31]~q ),
	.datad(!\M_rot_prestep2[23]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[7]~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[7]~27 .extended_lut = "off";
defparam \M_rot[7]~27 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[7]~27 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~27 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_mask[7]~q ),
	.datac(!\M_rot_pass1~q ),
	.datad(!\M_rot_sel_fill1~q ),
	.datae(!\M_rot[7]~27_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~27 .extended_lut = "off";
defparam \A_shift_rot_result~27 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~27 .shared_arith = "off";

dffeas \A_shift_rot_result[15] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~27_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_shift_rot_result[15]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[15] .is_wysiwyg = "true";
defparam \A_shift_rot_result[15] .power_up = "low";

dffeas \E_pc[13] (
	.clk(clk_clk),
	.d(\D_pc[13]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_pc[13]~q ),
	.prn(vcc));
defparam \E_pc[13] .is_wysiwyg = "true";
defparam \E_pc[13] .power_up = "low";

dffeas \E_pc[12] (
	.clk(clk_clk),
	.d(\D_pc[12]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_pc[12]~q ),
	.prn(vcc));
defparam \E_pc[12] .is_wysiwyg = "true";
defparam \E_pc[12] .power_up = "low";

dffeas \E_pc[11] (
	.clk(clk_clk),
	.d(\D_pc[11]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_pc[11]~q ),
	.prn(vcc));
defparam \E_pc[11] .is_wysiwyg = "true";
defparam \E_pc[11] .power_up = "low";

dffeas \E_pc[10] (
	.clk(clk_clk),
	.d(\D_pc[10]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_pc[10]~q ),
	.prn(vcc));
defparam \E_pc[10] .is_wysiwyg = "true";
defparam \E_pc[10] .power_up = "low";

cyclonev_lcell_comb \Add7~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_pc[10]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add7~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add7~45_sumout ),
	.cout(\Add7~46 ),
	.shareout());
defparam \Add7~45 .extended_lut = "off";
defparam \Add7~45 .lut_mask = 64'h00000000000000FF;
defparam \Add7~45 .shared_arith = "off";

cyclonev_lcell_comb \Add7~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_pc[11]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add7~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add7~49_sumout ),
	.cout(\Add7~50 ),
	.shareout());
defparam \Add7~49 .extended_lut = "off";
defparam \Add7~49 .lut_mask = 64'h00000000000000FF;
defparam \Add7~49 .shared_arith = "off";

cyclonev_lcell_comb \Add7~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_pc[12]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add7~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add7~53_sumout ),
	.cout(\Add7~54 ),
	.shareout());
defparam \Add7~53 .extended_lut = "off";
defparam \Add7~53 .lut_mask = 64'h00000000000000FF;
defparam \Add7~53 .shared_arith = "off";

cyclonev_lcell_comb \Add7~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_pc[13]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add7~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add7~41_sumout ),
	.cout(\Add7~42 ),
	.shareout());
defparam \Add7~41 .extended_lut = "off";
defparam \Add7~41 .lut_mask = 64'h00000000000000FF;
defparam \Add7~41 .shared_arith = "off";

dffeas \M_pc_plus_one[13] (
	.clk(clk_clk),
	.d(\Add7~41_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_pc_plus_one[13]~q ),
	.prn(vcc));
defparam \M_pc_plus_one[13] .is_wysiwyg = "true";
defparam \M_pc_plus_one[13] .power_up = "low";

dffeas \A_inst_result[15] (
	.clk(clk_clk),
	.d(\M_pc_plus_one[13]~q ),
	.asdata(\M_alu_result[15]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\A_inst_result[9]~0_combout ),
	.sload(!\M_exc_any~combout ),
	.ena(!\A_mem_stall~q ),
	.q(\A_inst_result[15]~q ),
	.prn(vcc));
defparam \A_inst_result[15] .is_wysiwyg = "true";
defparam \A_inst_result[15] .power_up = "low";

dffeas \A_mul_cell_p1[15] (
	.clk(clk_clk),
	.d(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[15]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_mul_cell_p1[15]~q ),
	.prn(vcc));
defparam \A_mul_cell_p1[15] .is_wysiwyg = "true";
defparam \A_mul_cell_p1[15] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[15]~29 (
	.dataa(!\A_slow_inst_result[15]~q ),
	.datab(!\A_shift_rot_result[15]~q ),
	.datac(!\A_inst_result[15]~q ),
	.datad(!\A_mul_cell_p1[15]~q ),
	.datae(!\A_wr_data_unfiltered[15]~0_combout ),
	.dataf(!\A_wr_data_unfiltered[15]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[15]~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[15]~29 .extended_lut = "off";
defparam \A_wr_data_unfiltered[15]~29 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_wr_data_unfiltered[15]~29 .shared_arith = "off";

dffeas \W_wr_data[15] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[15]~29_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[15]~q ),
	.prn(vcc));
defparam \W_wr_data[15] .is_wysiwyg = "true";
defparam \W_wr_data[15] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[15]~62 (
	.dataa(!\D_src2_reg[0]~7_combout ),
	.datab(!\D_src2_reg[0]~8_combout ),
	.datac(!\W_wr_data[15]~q ),
	.datad(!\A_wr_data_unfiltered[15]~29_combout ),
	.datae(!\M_alu_result[15]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[15]~62_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[15]~62 .extended_lut = "off";
defparam \D_src2_reg[15]~62 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \D_src2_reg[15]~62 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[15]~63 (
	.dataa(!\D_src2_reg[0]~4_combout ),
	.datab(!\D_src2_reg[0]~5_combout ),
	.datac(!\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[15] ),
	.datad(!\E_alu_result[15]~combout ),
	.datae(!\D_src2_reg[15]~62_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[15]~63_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[15]~63 .extended_lut = "off";
defparam \D_src2_reg[15]~63 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \D_src2_reg[15]~63 .shared_arith = "off";

dffeas \E_src2[15] (
	.clk(clk_clk),
	.d(\D_iw[21]~q ),
	.asdata(\D_src2_reg[15]~63_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src2[5]~2_combout ),
	.sload(!\D_ctrl_src2_choose_imm~q ),
	.ena(!\A_mem_stall~q ),
	.q(\E_src2[15]~q ),
	.prn(vcc));
defparam \E_src2[15] .is_wysiwyg = "true";
defparam \E_src2[15] .power_up = "low";

cyclonev_lcell_comb \Add9~29 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[12]~q ),
	.datae(gnd),
	.dataf(!\E_src1[12]~q ),
	.datag(gnd),
	.cin(\Add9~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~29_sumout ),
	.cout(\Add9~30 ),
	.shareout());
defparam \Add9~29 .extended_lut = "off";
defparam \Add9~29 .lut_mask = 64'h0000FF00000055AA;
defparam \Add9~29 .shared_arith = "off";

cyclonev_lcell_comb \Add9~25 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[13]~q ),
	.datae(gnd),
	.dataf(!\E_src1[13]~q ),
	.datag(gnd),
	.cin(\Add9~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~25_sumout ),
	.cout(\Add9~26 ),
	.shareout());
defparam \Add9~25 .extended_lut = "off";
defparam \Add9~25 .lut_mask = 64'h0000FF00000055AA;
defparam \Add9~25 .shared_arith = "off";

cyclonev_lcell_comb \Add9~21 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[14]~q ),
	.datae(gnd),
	.dataf(!\E_src1[14]~q ),
	.datag(gnd),
	.cin(\Add9~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~21_sumout ),
	.cout(\Add9~22 ),
	.shareout());
defparam \Add9~21 .extended_lut = "off";
defparam \Add9~21 .lut_mask = 64'h0000FF00000055AA;
defparam \Add9~21 .shared_arith = "off";

cyclonev_lcell_comb \Add9~17 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[15]~q ),
	.datae(gnd),
	.dataf(!\E_src1[15]~q ),
	.datag(gnd),
	.cin(\Add9~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~17_sumout ),
	.cout(\Add9~18 ),
	.shareout());
defparam \Add9~17 .extended_lut = "off";
defparam \Add9~17 .lut_mask = 64'h0000FF00000055AA;
defparam \Add9~17 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result~20 (
	.dataa(!\E_src2[15]~q ),
	.datab(!\E_src1[15]~q ),
	.datac(!\E_logic_op[1]~q ),
	.datad(!\E_logic_op[0]~q ),
	.datae(!\E_ctrl_logic~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result~20 .extended_lut = "off";
defparam \E_alu_result~20 .lut_mask = 64'h6996FFFF6996FFFF;
defparam \E_alu_result~20 .shared_arith = "off";

dffeas \E_extra_pc[13] (
	.clk(clk_clk),
	.d(\Add1~5_sumout ),
	.asdata(\D_pc_plus_one[13]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_br_pred_not_taken~combout ),
	.ena(!\A_mem_stall~q ),
	.q(\E_extra_pc[13]~q ),
	.prn(vcc));
defparam \E_extra_pc[13] .is_wysiwyg = "true";
defparam \E_extra_pc[13] .power_up = "low";

cyclonev_lcell_comb \E_alu_result[15] (
	.dataa(!\Add9~17_sumout ),
	.datab(!\E_ctrl_retaddr~q ),
	.datac(!\E_alu_result~0_combout ),
	.datad(!\E_alu_result~20_combout ),
	.datae(!\E_extra_pc[13]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[15]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[15] .extended_lut = "off";
defparam \E_alu_result[15] .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \E_alu_result[15] .shared_arith = "off";

dffeas \M_alu_result[15] (
	.clk(clk_clk),
	.d(\E_alu_result[15]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_alu_result[15]~q ),
	.prn(vcc));
defparam \M_alu_result[15] .is_wysiwyg = "true";
defparam \M_alu_result[15] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[15]~27 (
	.dataa(!\M_alu_result[15]~q ),
	.datab(!\A_wr_data_unfiltered[15]~29_combout ),
	.datac(!\first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[15] ),
	.datad(!\W_wr_data[15]~q ),
	.datae(!\E_src1[26]~0_combout ),
	.dataf(!\E_src1[26]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[15]~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[15]~27 .extended_lut = "off";
defparam \D_src1_reg[15]~27 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[15]~27 .shared_arith = "off";

dffeas \E_src1[15] (
	.clk(clk_clk),
	.d(\D_src1_reg[15]~27_combout ),
	.asdata(\E_alu_result[15]~combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\Equal303~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(!\A_mem_stall~q ),
	.q(\E_src1[15]~q ),
	.prn(vcc));
defparam \E_src1[15] .is_wysiwyg = "true";
defparam \E_src1[15] .power_up = "low";

cyclonev_lcell_comb \E_rot_step1[15]~28 (
	.dataa(!\E_src1[15]~q ),
	.datab(!\E_src1[14]~q ),
	.datac(!\E_src1[13]~q ),
	.datad(!\E_src1[12]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add10~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[15]~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[15]~28 .extended_lut = "off";
defparam \E_rot_step1[15]~28 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[15]~28 .shared_arith = "off";

dffeas \M_rot_prestep2[19] (
	.clk(clk_clk),
	.d(\E_rot_step1[15]~28_combout ),
	.asdata(\E_rot_step1[19]~29_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add10~1_combout ),
	.ena(!\A_mem_stall~q ),
	.q(\M_rot_prestep2[19]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[19] .is_wysiwyg = "true";
defparam \M_rot_prestep2[19] .power_up = "low";

cyclonev_lcell_comb \M_rot[3]~22 (
	.dataa(!\M_rot_prestep2[19]~q ),
	.datab(!\M_rot_prestep2[11]~q ),
	.datac(!\M_rot_prestep2[3]~q ),
	.datad(!\M_rot_prestep2[27]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[3]~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[3]~22 .extended_lut = "off";
defparam \M_rot[3]~22 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[3]~22 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~22 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_mask[3]~q ),
	.datac(!\M_rot_pass2~q ),
	.datad(!\M_rot_sel_fill2~q ),
	.datae(!\M_rot[3]~22_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~22 .extended_lut = "off";
defparam \A_shift_rot_result~22 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~22 .shared_arith = "off";

dffeas \A_shift_rot_result[19] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~22_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_shift_rot_result[19]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[19] .is_wysiwyg = "true";
defparam \A_shift_rot_result[19] .power_up = "low";

cyclonev_lcell_comb \A_inst_result[26]~1 (
	.dataa(!\M_exc_any~combout ),
	.datab(!\M_ctrl_rd_ctl_reg~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_inst_result[26]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_inst_result[26]~1 .extended_lut = "off";
defparam \A_inst_result[26]~1 .lut_mask = 64'h7777777777777777;
defparam \A_inst_result[26]~1 .shared_arith = "off";

dffeas \A_inst_result[19] (
	.clk(clk_clk),
	.d(\M_alu_result[19]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\A_inst_result[26]~1_combout ),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_inst_result[19]~q ),
	.prn(vcc));
defparam \A_inst_result[19] .is_wysiwyg = "true";
defparam \A_inst_result[19] .power_up = "low";

cyclonev_lcell_comb \Add11~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[0]~q ),
	.datae(gnd),
	.dataf(!\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[16]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add11~57_sumout ),
	.cout(\Add11~58 ),
	.shareout());
defparam \Add11~57 .extended_lut = "off";
defparam \Add11~57 .lut_mask = 64'h0000FF00000000FF;
defparam \Add11~57 .shared_arith = "off";

cyclonev_lcell_comb \Add11~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[1]~q ),
	.datae(gnd),
	.dataf(!\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[17]~q ),
	.datag(gnd),
	.cin(\Add11~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add11~45_sumout ),
	.cout(\Add11~46 ),
	.shareout());
defparam \Add11~45 .extended_lut = "off";
defparam \Add11~45 .lut_mask = 64'h0000FF00000000FF;
defparam \Add11~45 .shared_arith = "off";

cyclonev_lcell_comb \Add11~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[2]~q ),
	.datae(gnd),
	.dataf(!\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[18]~q ),
	.datag(gnd),
	.cin(\Add11~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add11~53_sumout ),
	.cout(\Add11~54 ),
	.shareout());
defparam \Add11~53 .extended_lut = "off";
defparam \Add11~53 .lut_mask = 64'h0000FF00000000FF;
defparam \Add11~53 .shared_arith = "off";

cyclonev_lcell_comb \Add11~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[3]~q ),
	.datae(gnd),
	.dataf(!\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[19]~q ),
	.datag(gnd),
	.cin(\Add11~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add11~41_sumout ),
	.cout(\Add11~42 ),
	.shareout());
defparam \Add11~41 .extended_lut = "off";
defparam \Add11~41 .lut_mask = 64'h0000FF00000000FF;
defparam \Add11~41 .shared_arith = "off";

dffeas \A_mul_s1[3] (
	.clk(clk_clk),
	.d(\Add11~41_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_mul_s1[3]~q ),
	.prn(vcc));
defparam \A_mul_s1[3] .is_wysiwyg = "true";
defparam \A_mul_s1[3] .power_up = "low";

dffeas \A_mul_cell_p3[3] (
	.clk(clk_clk),
	.d(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p3|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[3]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_mul_cell_p3[3]~q ),
	.prn(vcc));
defparam \A_mul_cell_p3[3] .is_wysiwyg = "true";
defparam \A_mul_cell_p3[3] .power_up = "low";

dffeas \A_mul_s1[2] (
	.clk(clk_clk),
	.d(\Add11~53_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_mul_s1[2]~q ),
	.prn(vcc));
defparam \A_mul_s1[2] .is_wysiwyg = "true";
defparam \A_mul_s1[2] .power_up = "low";

dffeas \A_mul_cell_p3[2] (
	.clk(clk_clk),
	.d(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p3|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[2]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_mul_cell_p3[2]~q ),
	.prn(vcc));
defparam \A_mul_cell_p3[2] .is_wysiwyg = "true";
defparam \A_mul_cell_p3[2] .power_up = "low";

dffeas \A_mul_s1[1] (
	.clk(clk_clk),
	.d(\Add11~45_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_mul_s1[1]~q ),
	.prn(vcc));
defparam \A_mul_s1[1] .is_wysiwyg = "true";
defparam \A_mul_s1[1] .power_up = "low";

dffeas \A_mul_cell_p3[1] (
	.clk(clk_clk),
	.d(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p3|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[1]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_mul_cell_p3[1]~q ),
	.prn(vcc));
defparam \A_mul_cell_p3[1] .is_wysiwyg = "true";
defparam \A_mul_cell_p3[1] .power_up = "low";

dffeas \A_mul_s1[0] (
	.clk(clk_clk),
	.d(\Add11~57_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_mul_s1[0]~q ),
	.prn(vcc));
defparam \A_mul_s1[0] .is_wysiwyg = "true";
defparam \A_mul_s1[0] .power_up = "low";

dffeas \A_mul_cell_p3[0] (
	.clk(clk_clk),
	.d(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p3|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[0]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_mul_cell_p3[0]~q ),
	.prn(vcc));
defparam \A_mul_cell_p3[0] .is_wysiwyg = "true";
defparam \A_mul_cell_p3[0] .power_up = "low";

cyclonev_lcell_comb \Add12~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_mul_s1[0]~q ),
	.datae(gnd),
	.dataf(!\A_mul_cell_p3[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add12~57_sumout ),
	.cout(\Add12~58 ),
	.shareout());
defparam \Add12~57 .extended_lut = "off";
defparam \Add12~57 .lut_mask = 64'h0000FF00000000FF;
defparam \Add12~57 .shared_arith = "off";

cyclonev_lcell_comb \Add12~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_mul_s1[1]~q ),
	.datae(gnd),
	.dataf(!\A_mul_cell_p3[1]~q ),
	.datag(gnd),
	.cin(\Add12~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add12~45_sumout ),
	.cout(\Add12~46 ),
	.shareout());
defparam \Add12~45 .extended_lut = "off";
defparam \Add12~45 .lut_mask = 64'h0000FF00000000FF;
defparam \Add12~45 .shared_arith = "off";

cyclonev_lcell_comb \Add12~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_mul_s1[2]~q ),
	.datae(gnd),
	.dataf(!\A_mul_cell_p3[2]~q ),
	.datag(gnd),
	.cin(\Add12~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add12~53_sumout ),
	.cout(\Add12~54 ),
	.shareout());
defparam \Add12~53 .extended_lut = "off";
defparam \Add12~53 .lut_mask = 64'h0000FF00000000FF;
defparam \Add12~53 .shared_arith = "off";

cyclonev_lcell_comb \Add12~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_mul_s1[3]~q ),
	.datae(gnd),
	.dataf(!\A_mul_cell_p3[3]~q ),
	.datag(gnd),
	.cin(\Add12~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add12~41_sumout ),
	.cout(\Add12~42 ),
	.shareout());
defparam \Add12~41 .extended_lut = "off";
defparam \Add12~41 .lut_mask = 64'h0000FF00000000FF;
defparam \Add12~41 .shared_arith = "off";

cyclonev_lcell_comb \A_wr_data_unfiltered[19]~24 (
	.dataa(!\A_slow_inst_result[19]~q ),
	.datab(!\A_shift_rot_result[19]~q ),
	.datac(!\A_inst_result[19]~q ),
	.datad(!\Add12~41_sumout ),
	.datae(!\A_wr_data_unfiltered[15]~0_combout ),
	.dataf(!\A_wr_data_unfiltered[15]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[19]~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[19]~24 .extended_lut = "off";
defparam \A_wr_data_unfiltered[19]~24 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_wr_data_unfiltered[19]~24 .shared_arith = "off";

dffeas \W_wr_data[19] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[19]~24_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[19]~q ),
	.prn(vcc));
defparam \W_wr_data[19] .is_wysiwyg = "true";
defparam \W_wr_data[19] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[19]~55 (
	.dataa(!\D_src2_reg[0]~4_combout ),
	.datab(!\D_src2_reg[0]~7_combout ),
	.datac(!\D_src2_reg[0]~8_combout ),
	.datad(!\M_alu_result[19]~q ),
	.datae(!\A_wr_data_unfiltered[19]~24_combout ),
	.dataf(!\W_wr_data[19]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[19]~55_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[19]~55 .extended_lut = "off";
defparam \D_src2_reg[19]~55 .lut_mask = 64'hBEFFFFFFFFFFFFFF;
defparam \D_src2_reg[19]~55 .shared_arith = "off";

cyclonev_lcell_comb \Add9~13 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[16]~q ),
	.datae(gnd),
	.dataf(!\E_src1[16]~q ),
	.datag(gnd),
	.cin(\Add9~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~13_sumout ),
	.cout(\Add9~14 ),
	.shareout());
defparam \Add9~13 .extended_lut = "off";
defparam \Add9~13 .lut_mask = 64'h0000FF00000055AA;
defparam \Add9~13 .shared_arith = "off";

cyclonev_lcell_comb \Add9~117 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[17]~q ),
	.datae(gnd),
	.dataf(!\E_src1[17]~q ),
	.datag(gnd),
	.cin(\Add9~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~117_sumout ),
	.cout(\Add9~118 ),
	.shareout());
defparam \Add9~117 .extended_lut = "off";
defparam \Add9~117 .lut_mask = 64'h0000FF00000055AA;
defparam \Add9~117 .shared_arith = "off";

cyclonev_lcell_comb \Add9~125 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[18]~q ),
	.datae(gnd),
	.dataf(!\E_src1[18]~q ),
	.datag(gnd),
	.cin(\Add9~118 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~125_sumout ),
	.cout(\Add9~126 ),
	.shareout());
defparam \Add9~125 .extended_lut = "off";
defparam \Add9~125 .lut_mask = 64'h0000FF00000055AA;
defparam \Add9~125 .shared_arith = "off";

cyclonev_lcell_comb \Add9~113 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[19]~q ),
	.datae(gnd),
	.dataf(!\E_src1[19]~q ),
	.datag(gnd),
	.cin(\Add9~126 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~113_sumout ),
	.cout(\Add9~114 ),
	.shareout());
defparam \Add9~113 .extended_lut = "off";
defparam \Add9~113 .lut_mask = 64'h0000FF00000055AA;
defparam \Add9~113 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~0 (
	.dataa(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[5] ),
	.datab(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[4] ),
	.datac(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[3] ),
	.datad(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[2] ),
	.datae(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[1] ),
	.dataf(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[0] ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~0 .extended_lut = "off";
defparam \Equal0~0 .lut_mask = 64'hFFFFFFFFFF7FFFFF;
defparam \Equal0~0 .shared_arith = "off";

cyclonev_lcell_comb \F_ctrl_unsigned_lo_imm16~1 (
	.dataa(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[5] ),
	.datab(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[4] ),
	.datac(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[3] ),
	.datad(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[2] ),
	.datae(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[0] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ctrl_unsigned_lo_imm16~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ctrl_unsigned_lo_imm16~1 .extended_lut = "off";
defparam \F_ctrl_unsigned_lo_imm16~1 .lut_mask = 64'hFFFF6996FFFF6996;
defparam \F_ctrl_unsigned_lo_imm16~1 .shared_arith = "off";

cyclonev_lcell_comb \F_ctrl_unsigned_lo_imm16~0 (
	.dataa(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[11] ),
	.datab(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[12] ),
	.datac(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[13] ),
	.datad(!\Equal0~0_combout ),
	.datae(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[1] ),
	.dataf(!\F_ctrl_unsigned_lo_imm16~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ctrl_unsigned_lo_imm16~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ctrl_unsigned_lo_imm16~0 .extended_lut = "off";
defparam \F_ctrl_unsigned_lo_imm16~0 .lut_mask = 64'hFFFFFBFFFFFFFFFF;
defparam \F_ctrl_unsigned_lo_imm16~0 .shared_arith = "off";

dffeas D_ctrl_unsigned_lo_imm16(
	.clk(clk_clk),
	.d(\F_ctrl_unsigned_lo_imm16~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_ctrl_unsigned_lo_imm16~q ),
	.prn(vcc));
defparam D_ctrl_unsigned_lo_imm16.is_wysiwyg = "true";
defparam D_ctrl_unsigned_lo_imm16.power_up = "low";

cyclonev_lcell_comb \D_src2[19]~37 (
	.dataa(!\D_ctrl_hi_imm16~q ),
	.datab(!\D_iw[21]~q ),
	.datac(!\D_ctrl_unsigned_lo_imm16~q ),
	.datad(!\D_iw[9]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[19]~37_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[19]~37 .extended_lut = "off";
defparam \D_src2[19]~37 .lut_mask = 64'h7BFF7BFF7BFF7BFF;
defparam \D_src2[19]~37 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[19]~38 (
	.dataa(!\D_ctrl_src2_choose_imm~q ),
	.datab(!\E_logic_result[19]~10_combout ),
	.datac(!\E_ctrl_logic~q ),
	.datad(!\E_alu_result~0_combout ),
	.datae(!\Add9~113_sumout ),
	.dataf(!\D_src2[19]~37_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[19]~38_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[19]~38 .extended_lut = "off";
defparam \D_src2[19]~38 .lut_mask = 64'h27FFFFFFFFFFFFFF;
defparam \D_src2[19]~38 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[19]~20 (
	.dataa(!\D_src2_reg[0]~5_combout ),
	.datab(!\D_ctrl_src2_choose_imm~q ),
	.datac(!\D_src2_reg[19]~55_combout ),
	.datad(!\D_src2_reg[0]~4_combout ),
	.datae(!\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[19] ),
	.dataf(!\D_src2[19]~38_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[19]~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[19]~20 .extended_lut = "off";
defparam \D_src2[19]~20 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \D_src2[19]~20 .shared_arith = "off";

cyclonev_lcell_comb \E_src2[30]~1 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\D_ctrl_src2_choose_imm~q ),
	.datac(!\D_ctrl_shift_right_arith~0_combout ),
	.datad(!\D_ctrl_unsigned_lo_imm16~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_src2[30]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_src2[30]~1 .extended_lut = "off";
defparam \E_src2[30]~1 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \E_src2[30]~1 .shared_arith = "off";

dffeas \E_src2[19] (
	.clk(clk_clk),
	.d(\D_src2[19]~20_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src2[30]~1_combout ),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_src2[19]~q ),
	.prn(vcc));
defparam \E_src2[19] .is_wysiwyg = "true";
defparam \E_src2[19] .power_up = "low";

cyclonev_lcell_comb \E_logic_result[19]~10 (
	.dataa(!\E_src2[19]~q ),
	.datab(!\E_src1[19]~q ),
	.datac(!\E_logic_op[1]~q ),
	.datad(!\E_logic_op[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[19]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[19]~10 .extended_lut = "off";
defparam \E_logic_result[19]~10 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[19]~10 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[19] (
	.dataa(!\E_logic_result[19]~10_combout ),
	.datab(!\E_ctrl_logic~q ),
	.datac(!\E_alu_result~0_combout ),
	.datad(!\Add9~113_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[19]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[19] .extended_lut = "off";
defparam \E_alu_result[19] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \E_alu_result[19] .shared_arith = "off";

dffeas \M_alu_result[19] (
	.clk(clk_clk),
	.d(\E_alu_result[19]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_alu_result[19]~q ),
	.prn(vcc));
defparam \M_alu_result[19] .is_wysiwyg = "true";
defparam \M_alu_result[19] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[19]~21 (
	.dataa(!\M_alu_result[19]~q ),
	.datab(!\A_wr_data_unfiltered[19]~24_combout ),
	.datac(!\first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[19] ),
	.datad(!\W_wr_data[19]~q ),
	.datae(!\E_src1[26]~0_combout ),
	.dataf(!\E_src1[26]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[19]~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[19]~21 .extended_lut = "off";
defparam \D_src1_reg[19]~21 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[19]~21 .shared_arith = "off";

dffeas \E_src1[19] (
	.clk(clk_clk),
	.d(\D_src1_reg[19]~21_combout ),
	.asdata(\E_alu_result[19]~combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\Equal303~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(!\A_mem_stall~q ),
	.q(\E_src1[19]~q ),
	.prn(vcc));
defparam \E_src1[19] .is_wysiwyg = "true";
defparam \E_src1[19] .power_up = "low";

cyclonev_lcell_comb \E_rot_step1[21]~10 (
	.dataa(!\E_src1[21]~q ),
	.datab(!\E_src1[20]~q ),
	.datac(!\E_src1[19]~q ),
	.datad(!\E_src1[18]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add10~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[21]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[21]~10 .extended_lut = "off";
defparam \E_rot_step1[21]~10 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[21]~10 .shared_arith = "off";

cyclonev_lcell_comb \E_rot_step1[25]~11 (
	.dataa(!\E_src1[25]~q ),
	.datab(!\E_src1[24]~q ),
	.datac(!\E_src1[23]~q ),
	.datad(!\E_src1[22]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add10~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[25]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[25]~11 .extended_lut = "off";
defparam \E_rot_step1[25]~11 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[25]~11 .shared_arith = "off";

dffeas \M_rot_prestep2[25] (
	.clk(clk_clk),
	.d(\E_rot_step1[21]~10_combout ),
	.asdata(\E_rot_step1[25]~11_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add10~1_combout ),
	.ena(!\A_mem_stall~q ),
	.q(\M_rot_prestep2[25]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[25] .is_wysiwyg = "true";
defparam \M_rot_prestep2[25] .power_up = "low";

cyclonev_lcell_comb \M_rot[1]~19 (
	.dataa(!\M_rot_prestep2[9]~q ),
	.datab(!\M_rot_prestep2[1]~q ),
	.datac(!\M_rot_prestep2[25]~q ),
	.datad(!\M_rot_prestep2[17]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[1]~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[1]~19 .extended_lut = "off";
defparam \M_rot[1]~19 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[1]~19 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~19 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_mask[1]~q ),
	.datac(!\M_rot_pass1~q ),
	.datad(!\M_rot_sel_fill1~q ),
	.datae(!\M_rot[1]~19_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~19 .extended_lut = "off";
defparam \A_shift_rot_result~19 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~19 .shared_arith = "off";

dffeas \A_shift_rot_result[9] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~19_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_shift_rot_result[9]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[9] .is_wysiwyg = "true";
defparam \A_shift_rot_result[9] .power_up = "low";

dffeas \M_pc_plus_one[7] (
	.clk(clk_clk),
	.d(\Add7~33_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_pc_plus_one[7]~q ),
	.prn(vcc));
defparam \M_pc_plus_one[7] .is_wysiwyg = "true";
defparam \M_pc_plus_one[7] .power_up = "low";

dffeas \A_inst_result[9] (
	.clk(clk_clk),
	.d(\M_pc_plus_one[7]~q ),
	.asdata(\M_alu_result[9]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\A_inst_result[9]~0_combout ),
	.sload(!\M_exc_any~combout ),
	.ena(!\A_mem_stall~q ),
	.q(\A_inst_result[9]~q ),
	.prn(vcc));
defparam \A_inst_result[9] .is_wysiwyg = "true";
defparam \A_inst_result[9] .power_up = "low";

dffeas \A_mul_cell_p1[9] (
	.clk(clk_clk),
	.d(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[9]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_mul_cell_p1[9]~q ),
	.prn(vcc));
defparam \A_mul_cell_p1[9] .is_wysiwyg = "true";
defparam \A_mul_cell_p1[9] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[9]~21 (
	.dataa(!\A_slow_inst_result[9]~q ),
	.datab(!\A_shift_rot_result[9]~q ),
	.datac(!\A_inst_result[9]~q ),
	.datad(!\A_mul_cell_p1[9]~q ),
	.datae(!\A_wr_data_unfiltered[15]~0_combout ),
	.dataf(!\A_wr_data_unfiltered[15]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[9]~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[9]~21 .extended_lut = "off";
defparam \A_wr_data_unfiltered[9]~21 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_wr_data_unfiltered[9]~21 .shared_arith = "off";

dffeas \W_wr_data[9] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[9]~21_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[9]~q ),
	.prn(vcc));
defparam \W_wr_data[9] .is_wysiwyg = "true";
defparam \W_wr_data[9] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[9]~50 (
	.dataa(!\D_src2_reg[0]~7_combout ),
	.datab(!\D_src2_reg[0]~8_combout ),
	.datac(!\W_wr_data[9]~q ),
	.datad(!\A_wr_data_unfiltered[9]~21_combout ),
	.datae(!\M_alu_result[9]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[9]~50_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[9]~50 .extended_lut = "off";
defparam \D_src2_reg[9]~50 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \D_src2_reg[9]~50 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[9]~51 (
	.dataa(!\D_src2_reg[0]~4_combout ),
	.datab(!\D_src2_reg[0]~5_combout ),
	.datac(!\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[9] ),
	.datad(!\E_alu_result[9]~combout ),
	.datae(!\D_src2_reg[9]~50_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[9]~51_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[9]~51 .extended_lut = "off";
defparam \D_src2_reg[9]~51 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \D_src2_reg[9]~51 .shared_arith = "off";

dffeas \E_src2[9] (
	.clk(clk_clk),
	.d(\D_iw[15]~q ),
	.asdata(\D_src2_reg[9]~51_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src2[5]~2_combout ),
	.sload(!\D_ctrl_src2_choose_imm~q ),
	.ena(!\A_mem_stall~q ),
	.q(\E_src2[9]~q ),
	.prn(vcc));
defparam \E_src2[9] .is_wysiwyg = "true";
defparam \E_src2[9] .power_up = "low";

cyclonev_lcell_comb \E_alu_result~16 (
	.dataa(!\E_src2[9]~q ),
	.datab(!\E_src1[9]~q ),
	.datac(!\E_logic_op[1]~q ),
	.datad(!\E_logic_op[0]~q ),
	.datae(!\E_ctrl_logic~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result~16 .extended_lut = "off";
defparam \E_alu_result~16 .lut_mask = 64'h6996FFFF6996FFFF;
defparam \E_alu_result~16 .shared_arith = "off";

dffeas \D_pc_plus_one[7] (
	.clk(clk_clk),
	.d(\Add3~29_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_pc_plus_one[7]~q ),
	.prn(vcc));
defparam \D_pc_plus_one[7] .is_wysiwyg = "true";
defparam \D_pc_plus_one[7] .power_up = "low";

dffeas \E_extra_pc[7] (
	.clk(clk_clk),
	.d(\D_br_taken_waddr_partial[7]~q ),
	.asdata(\D_pc_plus_one[7]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_br_pred_not_taken~combout ),
	.ena(!\A_mem_stall~q ),
	.q(\E_extra_pc[7]~q ),
	.prn(vcc));
defparam \E_extra_pc[7] .is_wysiwyg = "true";
defparam \E_extra_pc[7] .power_up = "low";

cyclonev_lcell_comb \E_alu_result[9] (
	.dataa(!\Add9~41_sumout ),
	.datab(!\E_ctrl_retaddr~q ),
	.datac(!\E_alu_result~0_combout ),
	.datad(!\E_alu_result~16_combout ),
	.datae(!\E_extra_pc[7]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[9]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[9] .extended_lut = "off";
defparam \E_alu_result[9] .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \E_alu_result[9] .shared_arith = "off";

dffeas \M_alu_result[9] (
	.clk(clk_clk),
	.d(\E_alu_result[9]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_alu_result[9]~q ),
	.prn(vcc));
defparam \M_alu_result[9] .is_wysiwyg = "true";
defparam \M_alu_result[9] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[9]~15 (
	.dataa(!\M_alu_result[9]~q ),
	.datab(!\A_wr_data_unfiltered[9]~21_combout ),
	.datac(!\first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[9] ),
	.datad(!\W_wr_data[9]~q ),
	.datae(!\E_src1[26]~0_combout ),
	.dataf(!\E_src1[26]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[9]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[9]~15 .extended_lut = "off";
defparam \D_src1_reg[9]~15 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[9]~15 .shared_arith = "off";

dffeas \E_src1[9] (
	.clk(clk_clk),
	.d(\D_src1_reg[9]~15_combout ),
	.asdata(\E_alu_result[9]~combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\Equal303~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(!\A_mem_stall~q ),
	.q(\E_src1[9]~q ),
	.prn(vcc));
defparam \E_src1[9] .is_wysiwyg = "true";
defparam \E_src1[9] .power_up = "low";

cyclonev_lcell_comb \E_rot_step1[9]~15 (
	.dataa(!\E_src1[9]~q ),
	.datab(!\E_src1[8]~q ),
	.datac(!\E_src1[7]~q ),
	.datad(!\E_src1[6]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add10~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[9]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[9]~15 .extended_lut = "off";
defparam \E_rot_step1[9]~15 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[9]~15 .shared_arith = "off";

dffeas \M_rot_prestep2[13] (
	.clk(clk_clk),
	.d(\E_rot_step1[9]~15_combout ),
	.asdata(\E_rot_step1[13]~12_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add10~1_combout ),
	.ena(!\A_mem_stall~q ),
	.q(\M_rot_prestep2[13]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[13] .is_wysiwyg = "true";
defparam \M_rot_prestep2[13] .power_up = "low";

dffeas \M_rot_prestep2[29] (
	.clk(clk_clk),
	.d(\E_rot_step1[25]~11_combout ),
	.asdata(\E_rot_step1[29]~8_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add10~1_combout ),
	.ena(!\A_mem_stall~q ),
	.q(\M_rot_prestep2[29]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[29] .is_wysiwyg = "true";
defparam \M_rot_prestep2[29] .power_up = "low";

cyclonev_lcell_comb \M_rot[5]~29 (
	.dataa(!\M_rot_prestep2[13]~q ),
	.datab(!\M_rot_prestep2[5]~q ),
	.datac(!\M_rot_prestep2[29]~q ),
	.datad(!\M_rot_prestep2[21]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[5]~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[5]~29 .extended_lut = "off";
defparam \M_rot[5]~29 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[5]~29 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~29 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_mask[5]~q ),
	.datac(!\M_rot_pass1~q ),
	.datad(!\M_rot_sel_fill1~q ),
	.datae(!\M_rot[5]~29_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~29 .extended_lut = "off";
defparam \A_shift_rot_result~29 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~29 .shared_arith = "off";

dffeas \A_shift_rot_result[13] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~29_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_shift_rot_result[13]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[13] .is_wysiwyg = "true";
defparam \A_shift_rot_result[13] .power_up = "low";

dffeas \M_pc_plus_one[11] (
	.clk(clk_clk),
	.d(\Add7~49_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_pc_plus_one[11]~q ),
	.prn(vcc));
defparam \M_pc_plus_one[11] .is_wysiwyg = "true";
defparam \M_pc_plus_one[11] .power_up = "low";

dffeas \A_inst_result[13] (
	.clk(clk_clk),
	.d(\M_pc_plus_one[11]~q ),
	.asdata(\M_alu_result[13]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\A_inst_result[9]~0_combout ),
	.sload(!\M_exc_any~combout ),
	.ena(!\A_mem_stall~q ),
	.q(\A_inst_result[13]~q ),
	.prn(vcc));
defparam \A_inst_result[13] .is_wysiwyg = "true";
defparam \A_inst_result[13] .power_up = "low";

dffeas \A_mul_cell_p1[13] (
	.clk(clk_clk),
	.d(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[13]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_mul_cell_p1[13]~q ),
	.prn(vcc));
defparam \A_mul_cell_p1[13] .is_wysiwyg = "true";
defparam \A_mul_cell_p1[13] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[13]~31 (
	.dataa(!\A_slow_inst_result[13]~q ),
	.datab(!\A_shift_rot_result[13]~q ),
	.datac(!\A_inst_result[13]~q ),
	.datad(!\A_mul_cell_p1[13]~q ),
	.datae(!\A_wr_data_unfiltered[15]~0_combout ),
	.dataf(!\A_wr_data_unfiltered[15]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[13]~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[13]~31 .extended_lut = "off";
defparam \A_wr_data_unfiltered[13]~31 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_wr_data_unfiltered[13]~31 .shared_arith = "off";

dffeas \W_wr_data[13] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[13]~31_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[13]~q ),
	.prn(vcc));
defparam \W_wr_data[13] .is_wysiwyg = "true";
defparam \W_wr_data[13] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[13]~66 (
	.dataa(!\D_src2_reg[0]~7_combout ),
	.datab(!\D_src2_reg[0]~8_combout ),
	.datac(!\W_wr_data[13]~q ),
	.datad(!\A_wr_data_unfiltered[13]~31_combout ),
	.datae(!\M_alu_result[13]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[13]~66_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[13]~66 .extended_lut = "off";
defparam \D_src2_reg[13]~66 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \D_src2_reg[13]~66 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[13]~67 (
	.dataa(!\D_src2_reg[0]~4_combout ),
	.datab(!\D_src2_reg[0]~5_combout ),
	.datac(!\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[13] ),
	.datad(!\E_alu_result[13]~combout ),
	.datae(!\D_src2_reg[13]~66_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[13]~67_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[13]~67 .extended_lut = "off";
defparam \D_src2_reg[13]~67 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \D_src2_reg[13]~67 .shared_arith = "off";

dffeas \E_src2[13] (
	.clk(clk_clk),
	.d(\D_iw[19]~q ),
	.asdata(\D_src2_reg[13]~67_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src2[5]~2_combout ),
	.sload(!\D_ctrl_src2_choose_imm~q ),
	.ena(!\A_mem_stall~q ),
	.q(\E_src2[13]~q ),
	.prn(vcc));
defparam \E_src2[13] .is_wysiwyg = "true";
defparam \E_src2[13] .power_up = "low";

cyclonev_lcell_comb \E_alu_result~22 (
	.dataa(!\E_src2[13]~q ),
	.datab(!\E_src1[13]~q ),
	.datac(!\E_logic_op[1]~q ),
	.datad(!\E_logic_op[0]~q ),
	.datae(!\E_ctrl_logic~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result~22 .extended_lut = "off";
defparam \E_alu_result~22 .lut_mask = 64'h6996FFFF6996FFFF;
defparam \E_alu_result~22 .shared_arith = "off";

dffeas \E_extra_pc[11] (
	.clk(clk_clk),
	.d(\Add1~13_sumout ),
	.asdata(\D_pc_plus_one[11]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_br_pred_not_taken~combout ),
	.ena(!\A_mem_stall~q ),
	.q(\E_extra_pc[11]~q ),
	.prn(vcc));
defparam \E_extra_pc[11] .is_wysiwyg = "true";
defparam \E_extra_pc[11] .power_up = "low";

cyclonev_lcell_comb \E_alu_result[13] (
	.dataa(!\Add9~25_sumout ),
	.datab(!\E_ctrl_retaddr~q ),
	.datac(!\E_alu_result~0_combout ),
	.datad(!\E_alu_result~22_combout ),
	.datae(!\E_extra_pc[11]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[13]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[13] .extended_lut = "off";
defparam \E_alu_result[13] .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \E_alu_result[13] .shared_arith = "off";

dffeas \M_alu_result[13] (
	.clk(clk_clk),
	.d(\E_alu_result[13]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_alu_result[13]~q ),
	.prn(vcc));
defparam \M_alu_result[13] .is_wysiwyg = "true";
defparam \M_alu_result[13] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[13]~29 (
	.dataa(!\M_alu_result[13]~q ),
	.datab(!\A_wr_data_unfiltered[13]~31_combout ),
	.datac(!\first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[13] ),
	.datad(!\W_wr_data[13]~q ),
	.datae(!\E_src1[26]~0_combout ),
	.dataf(!\E_src1[26]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[13]~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[13]~29 .extended_lut = "off";
defparam \D_src1_reg[13]~29 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[13]~29 .shared_arith = "off";

dffeas \E_src1[13] (
	.clk(clk_clk),
	.d(\D_src1_reg[13]~29_combout ),
	.asdata(\E_alu_result[13]~combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\Equal303~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(!\A_mem_stall~q ),
	.q(\E_src1[13]~q ),
	.prn(vcc));
defparam \E_src1[13] .is_wysiwyg = "true";
defparam \E_src1[13] .power_up = "low";

cyclonev_lcell_comb \E_rot_step1[13]~12 (
	.dataa(!\E_src1[13]~q ),
	.datab(!\E_src1[12]~q ),
	.datac(!\E_src1[11]~q ),
	.datad(!\E_src1[10]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add10~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[13]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[13]~12 .extended_lut = "off";
defparam \E_rot_step1[13]~12 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[13]~12 .shared_arith = "off";

dffeas \M_rot_prestep2[17] (
	.clk(clk_clk),
	.d(\E_rot_step1[13]~12_combout ),
	.asdata(\E_rot_step1[17]~13_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add10~1_combout ),
	.ena(!\A_mem_stall~q ),
	.q(\M_rot_prestep2[17]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[17] .is_wysiwyg = "true";
defparam \M_rot_prestep2[17] .power_up = "low";

cyclonev_lcell_comb \M_rot[1]~23 (
	.dataa(!\M_rot_prestep2[17]~q ),
	.datab(!\M_rot_prestep2[9]~q ),
	.datac(!\M_rot_prestep2[1]~q ),
	.datad(!\M_rot_prestep2[25]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[1]~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[1]~23 .extended_lut = "off";
defparam \M_rot[1]~23 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[1]~23 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~23 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_mask[1]~q ),
	.datac(!\M_rot_pass2~q ),
	.datad(!\M_rot_sel_fill2~q ),
	.datae(!\M_rot[1]~23_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~23 .extended_lut = "off";
defparam \A_shift_rot_result~23 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~23 .shared_arith = "off";

dffeas \A_shift_rot_result[17] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~23_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_shift_rot_result[17]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[17] .is_wysiwyg = "true";
defparam \A_shift_rot_result[17] .power_up = "low";

dffeas \A_inst_result[17] (
	.clk(clk_clk),
	.d(\M_alu_result[17]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\A_inst_result[26]~1_combout ),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_inst_result[17]~q ),
	.prn(vcc));
defparam \A_inst_result[17] .is_wysiwyg = "true";
defparam \A_inst_result[17] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[17]~25 (
	.dataa(!\A_slow_inst_result[17]~q ),
	.datab(!\A_shift_rot_result[17]~q ),
	.datac(!\A_inst_result[17]~q ),
	.datad(!\Add12~45_sumout ),
	.datae(!\A_wr_data_unfiltered[15]~0_combout ),
	.dataf(!\A_wr_data_unfiltered[15]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[17]~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[17]~25 .extended_lut = "off";
defparam \A_wr_data_unfiltered[17]~25 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_wr_data_unfiltered[17]~25 .shared_arith = "off";

dffeas \W_wr_data[17] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[17]~25_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[17]~q ),
	.prn(vcc));
defparam \W_wr_data[17] .is_wysiwyg = "true";
defparam \W_wr_data[17] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[17]~56 (
	.dataa(!\D_src2_reg[0]~4_combout ),
	.datab(!\D_src2_reg[0]~7_combout ),
	.datac(!\D_src2_reg[0]~8_combout ),
	.datad(!\M_alu_result[17]~q ),
	.datae(!\A_wr_data_unfiltered[17]~25_combout ),
	.dataf(!\W_wr_data[17]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[17]~56_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[17]~56 .extended_lut = "off";
defparam \D_src2_reg[17]~56 .lut_mask = 64'hBEFFFFFFFFFFFFFF;
defparam \D_src2_reg[17]~56 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[17]~33 (
	.dataa(!\D_ctrl_hi_imm16~q ),
	.datab(!\D_iw[21]~q ),
	.datac(!\D_ctrl_unsigned_lo_imm16~q ),
	.datad(!\D_iw[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[17]~33_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[17]~33 .extended_lut = "off";
defparam \D_src2[17]~33 .lut_mask = 64'h7BFF7BFF7BFF7BFF;
defparam \D_src2[17]~33 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[17]~34 (
	.dataa(!\D_ctrl_src2_choose_imm~q ),
	.datab(!\E_logic_result[17]~4_combout ),
	.datac(!\E_ctrl_logic~q ),
	.datad(!\E_alu_result~0_combout ),
	.datae(!\Add9~117_sumout ),
	.dataf(!\D_src2[17]~33_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[17]~34_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[17]~34 .extended_lut = "off";
defparam \D_src2[17]~34 .lut_mask = 64'h27FFFFFFFFFFFFFF;
defparam \D_src2[17]~34 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[17]~21 (
	.dataa(!\D_src2_reg[0]~5_combout ),
	.datab(!\D_ctrl_src2_choose_imm~q ),
	.datac(!\D_src2_reg[17]~56_combout ),
	.datad(!\D_src2_reg[0]~4_combout ),
	.datae(!\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[17] ),
	.dataf(!\D_src2[17]~34_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[17]~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[17]~21 .extended_lut = "off";
defparam \D_src2[17]~21 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \D_src2[17]~21 .shared_arith = "off";

dffeas \E_src2[17] (
	.clk(clk_clk),
	.d(\D_src2[17]~21_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src2[30]~1_combout ),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_src2[17]~q ),
	.prn(vcc));
defparam \E_src2[17] .is_wysiwyg = "true";
defparam \E_src2[17] .power_up = "low";

cyclonev_lcell_comb \E_logic_result[17]~4 (
	.dataa(!\E_src2[17]~q ),
	.datab(!\E_src1[17]~q ),
	.datac(!\E_logic_op[1]~q ),
	.datad(!\E_logic_op[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[17]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[17]~4 .extended_lut = "off";
defparam \E_logic_result[17]~4 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[17]~4 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[17] (
	.dataa(!\E_logic_result[17]~4_combout ),
	.datab(!\E_ctrl_logic~q ),
	.datac(!\E_alu_result~0_combout ),
	.datad(!\Add9~117_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[17]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[17] .extended_lut = "off";
defparam \E_alu_result[17] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \E_alu_result[17] .shared_arith = "off";

dffeas \M_alu_result[17] (
	.clk(clk_clk),
	.d(\E_alu_result[17]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_alu_result[17]~q ),
	.prn(vcc));
defparam \M_alu_result[17] .is_wysiwyg = "true";
defparam \M_alu_result[17] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[17]~22 (
	.dataa(!\M_alu_result[17]~q ),
	.datab(!\A_wr_data_unfiltered[17]~25_combout ),
	.datac(!\first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[17] ),
	.datad(!\W_wr_data[17]~q ),
	.datae(!\E_src1[26]~0_combout ),
	.dataf(!\E_src1[26]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[17]~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[17]~22 .extended_lut = "off";
defparam \D_src1_reg[17]~22 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[17]~22 .shared_arith = "off";

dffeas \E_src1[17] (
	.clk(clk_clk),
	.d(\D_src1_reg[17]~22_combout ),
	.asdata(\E_alu_result[17]~combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\Equal303~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(!\A_mem_stall~q ),
	.q(\E_src1[17]~q ),
	.prn(vcc));
defparam \E_src1[17] .is_wysiwyg = "true";
defparam \E_src1[17] .power_up = "low";

cyclonev_lcell_comb \E_rot_step1[17]~13 (
	.dataa(!\E_src1[17]~q ),
	.datab(!\E_src1[16]~q ),
	.datac(!\E_src1[15]~q ),
	.datad(!\E_src1[14]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add10~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[17]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[17]~13 .extended_lut = "off";
defparam \E_rot_step1[17]~13 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[17]~13 .shared_arith = "off";

dffeas \M_rot_prestep2[21] (
	.clk(clk_clk),
	.d(\E_rot_step1[17]~13_combout ),
	.asdata(\E_rot_step1[21]~10_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add10~1_combout ),
	.ena(!\A_mem_stall~q ),
	.q(\M_rot_prestep2[21]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[21] .is_wysiwyg = "true";
defparam \M_rot_prestep2[21] .power_up = "low";

cyclonev_lcell_comb \M_rot[5]~13 (
	.dataa(!\M_rot_prestep2[21]~q ),
	.datab(!\M_rot_prestep2[13]~q ),
	.datac(!\M_rot_prestep2[5]~q ),
	.datad(!\M_rot_prestep2[29]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[5]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[5]~13 .extended_lut = "off";
defparam \M_rot[5]~13 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[5]~13 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~13 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_mask[5]~q ),
	.datac(!\M_rot_pass2~q ),
	.datad(!\M_rot_sel_fill2~q ),
	.datae(!\M_rot[5]~13_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~13 .extended_lut = "off";
defparam \A_shift_rot_result~13 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~13 .shared_arith = "off";

dffeas \A_shift_rot_result[21] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~13_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_shift_rot_result[21]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[21] .is_wysiwyg = "true";
defparam \A_shift_rot_result[21] .power_up = "low";

dffeas \A_inst_result[21] (
	.clk(clk_clk),
	.d(\M_alu_result[21]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\A_inst_result[26]~1_combout ),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_inst_result[21]~q ),
	.prn(vcc));
defparam \A_inst_result[21] .is_wysiwyg = "true";
defparam \A_inst_result[21] .power_up = "low";

cyclonev_lcell_comb \Add11~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[4]~q ),
	.datae(gnd),
	.dataf(!\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[20]~q ),
	.datag(gnd),
	.cin(\Add11~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add11~37_sumout ),
	.cout(\Add11~38 ),
	.shareout());
defparam \Add11~37 .extended_lut = "off";
defparam \Add11~37 .lut_mask = 64'h0000FF00000000FF;
defparam \Add11~37 .shared_arith = "off";

cyclonev_lcell_comb \Add11~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[5]~q ),
	.datae(gnd),
	.dataf(!\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[21]~q ),
	.datag(gnd),
	.cin(\Add11~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add11~21_sumout ),
	.cout(\Add11~22 ),
	.shareout());
defparam \Add11~21 .extended_lut = "off";
defparam \Add11~21 .lut_mask = 64'h0000FF00000000FF;
defparam \Add11~21 .shared_arith = "off";

dffeas \A_mul_s1[5] (
	.clk(clk_clk),
	.d(\Add11~21_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_mul_s1[5]~q ),
	.prn(vcc));
defparam \A_mul_s1[5] .is_wysiwyg = "true";
defparam \A_mul_s1[5] .power_up = "low";

dffeas \A_mul_cell_p3[5] (
	.clk(clk_clk),
	.d(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p3|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[5]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_mul_cell_p3[5]~q ),
	.prn(vcc));
defparam \A_mul_cell_p3[5] .is_wysiwyg = "true";
defparam \A_mul_cell_p3[5] .power_up = "low";

dffeas \A_mul_s1[4] (
	.clk(clk_clk),
	.d(\Add11~37_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_mul_s1[4]~q ),
	.prn(vcc));
defparam \A_mul_s1[4] .is_wysiwyg = "true";
defparam \A_mul_s1[4] .power_up = "low";

dffeas \A_mul_cell_p3[4] (
	.clk(clk_clk),
	.d(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p3|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[4]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_mul_cell_p3[4]~q ),
	.prn(vcc));
defparam \A_mul_cell_p3[4] .is_wysiwyg = "true";
defparam \A_mul_cell_p3[4] .power_up = "low";

cyclonev_lcell_comb \Add12~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_mul_s1[4]~q ),
	.datae(gnd),
	.dataf(!\A_mul_cell_p3[4]~q ),
	.datag(gnd),
	.cin(\Add12~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add12~37_sumout ),
	.cout(\Add12~38 ),
	.shareout());
defparam \Add12~37 .extended_lut = "off";
defparam \Add12~37 .lut_mask = 64'h0000FF00000000FF;
defparam \Add12~37 .shared_arith = "off";

cyclonev_lcell_comb \Add12~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_mul_s1[5]~q ),
	.datae(gnd),
	.dataf(!\A_mul_cell_p3[5]~q ),
	.datag(gnd),
	.cin(\Add12~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add12~21_sumout ),
	.cout(\Add12~22 ),
	.shareout());
defparam \Add12~21 .extended_lut = "off";
defparam \Add12~21 .lut_mask = 64'h0000FF00000000FF;
defparam \Add12~21 .shared_arith = "off";

cyclonev_lcell_comb \A_wr_data_unfiltered[21]~15 (
	.dataa(!\A_slow_inst_result[21]~q ),
	.datab(!\A_shift_rot_result[21]~q ),
	.datac(!\A_inst_result[21]~q ),
	.datad(!\Add12~21_sumout ),
	.datae(!\A_wr_data_unfiltered[15]~0_combout ),
	.dataf(!\A_wr_data_unfiltered[15]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[21]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[21]~15 .extended_lut = "off";
defparam \A_wr_data_unfiltered[21]~15 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_wr_data_unfiltered[21]~15 .shared_arith = "off";

dffeas \W_wr_data[21] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[21]~15_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[21]~q ),
	.prn(vcc));
defparam \W_wr_data[21] .is_wysiwyg = "true";
defparam \W_wr_data[21] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[21]~37 (
	.dataa(!\D_src2_reg[0]~4_combout ),
	.datab(!\D_src2_reg[0]~7_combout ),
	.datac(!\D_src2_reg[0]~8_combout ),
	.datad(!\M_alu_result[21]~q ),
	.datae(!\A_wr_data_unfiltered[21]~15_combout ),
	.dataf(!\W_wr_data[21]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[21]~37_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[21]~37 .extended_lut = "off";
defparam \D_src2_reg[21]~37 .lut_mask = 64'hBEFFFFFFFFFFFFFF;
defparam \D_src2_reg[21]~37 .shared_arith = "off";

cyclonev_lcell_comb \Add9~109 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[20]~q ),
	.datae(gnd),
	.dataf(!\E_src1[20]~q ),
	.datag(gnd),
	.cin(\Add9~114 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~109_sumout ),
	.cout(\Add9~110 ),
	.shareout());
defparam \Add9~109 .extended_lut = "off";
defparam \Add9~109 .lut_mask = 64'h0000FF00000055AA;
defparam \Add9~109 .shared_arith = "off";

cyclonev_lcell_comb \Add9~93 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[21]~q ),
	.datae(gnd),
	.dataf(!\E_src1[21]~q ),
	.datag(gnd),
	.cin(\Add9~110 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~93_sumout ),
	.cout(\Add9~94 ),
	.shareout());
defparam \Add9~93 .extended_lut = "off";
defparam \Add9~93 .lut_mask = 64'h0000FF00000055AA;
defparam \Add9~93 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[21]~29 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\D_ctrl_hi_imm16~q ),
	.datac(!\D_iw[21]~q ),
	.datad(!\D_ctrl_unsigned_lo_imm16~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[21]~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[21]~29 .extended_lut = "off";
defparam \D_src2[21]~29 .lut_mask = 64'h7FDF7FDF7FDF7FDF;
defparam \D_src2[21]~29 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[21]~30 (
	.dataa(!\D_ctrl_src2_choose_imm~q ),
	.datab(!\E_logic_result[21]~8_combout ),
	.datac(!\E_ctrl_logic~q ),
	.datad(!\E_alu_result~0_combout ),
	.datae(!\Add9~93_sumout ),
	.dataf(!\D_src2[21]~29_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[21]~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[21]~30 .extended_lut = "off";
defparam \D_src2[21]~30 .lut_mask = 64'h27FFFFFFFFFFFFFF;
defparam \D_src2[21]~30 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[21]~11 (
	.dataa(!\D_src2_reg[0]~5_combout ),
	.datab(!\D_ctrl_src2_choose_imm~q ),
	.datac(!\D_src2_reg[21]~37_combout ),
	.datad(!\D_src2_reg[0]~4_combout ),
	.datae(!\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[21] ),
	.dataf(!\D_src2[21]~30_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[21]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[21]~11 .extended_lut = "off";
defparam \D_src2[21]~11 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \D_src2[21]~11 .shared_arith = "off";

dffeas \E_src2[21] (
	.clk(clk_clk),
	.d(\D_src2[21]~11_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src2[30]~1_combout ),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_src2[21]~q ),
	.prn(vcc));
defparam \E_src2[21] .is_wysiwyg = "true";
defparam \E_src2[21] .power_up = "low";

cyclonev_lcell_comb \E_logic_result[21]~8 (
	.dataa(!\E_src2[21]~q ),
	.datab(!\E_src1[21]~q ),
	.datac(!\E_logic_op[1]~q ),
	.datad(!\E_logic_op[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[21]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[21]~8 .extended_lut = "off";
defparam \E_logic_result[21]~8 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[21]~8 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[21] (
	.dataa(!\E_logic_result[21]~8_combout ),
	.datab(!\E_ctrl_logic~q ),
	.datac(!\E_alu_result~0_combout ),
	.datad(!\Add9~93_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[21]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[21] .extended_lut = "off";
defparam \E_alu_result[21] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \E_alu_result[21] .shared_arith = "off";

dffeas \M_alu_result[21] (
	.clk(clk_clk),
	.d(\E_alu_result[21]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_alu_result[21]~q ),
	.prn(vcc));
defparam \M_alu_result[21] .is_wysiwyg = "true";
defparam \M_alu_result[21] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[21]~9 (
	.dataa(!\M_alu_result[21]~q ),
	.datab(!\A_wr_data_unfiltered[21]~15_combout ),
	.datac(!\first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[21] ),
	.datad(!\W_wr_data[21]~q ),
	.datae(!\E_src1[26]~0_combout ),
	.dataf(!\E_src1[26]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[21]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[21]~9 .extended_lut = "off";
defparam \D_src1_reg[21]~9 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[21]~9 .shared_arith = "off";

dffeas \E_src1[21] (
	.clk(clk_clk),
	.d(\D_src1_reg[21]~9_combout ),
	.asdata(\E_alu_result[21]~combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\Equal303~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(!\A_mem_stall~q ),
	.q(\E_src1[21]~q ),
	.prn(vcc));
defparam \E_src1[21] .is_wysiwyg = "true";
defparam \E_src1[21] .power_up = "low";

cyclonev_lcell_comb \E_rot_step1[24]~3 (
	.dataa(!\E_src1[24]~q ),
	.datab(!\E_src1[23]~q ),
	.datac(!\E_src1[22]~q ),
	.datad(!\E_src1[21]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add10~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[24]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[24]~3 .extended_lut = "off";
defparam \E_rot_step1[24]~3 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[24]~3 .shared_arith = "off";

dffeas \M_rot_prestep2[28] (
	.clk(clk_clk),
	.d(\E_rot_step1[24]~3_combout ),
	.asdata(\E_rot_step1[28]~0_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add10~1_combout ),
	.ena(!\A_mem_stall~q ),
	.q(\M_rot_prestep2[28]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[28] .is_wysiwyg = "true";
defparam \M_rot_prestep2[28] .power_up = "low";

cyclonev_lcell_comb \M_rot[4]~28 (
	.dataa(!\M_rot_prestep2[12]~q ),
	.datab(!\M_rot_prestep2[4]~q ),
	.datac(!\M_rot_prestep2[28]~q ),
	.datad(!\M_rot_prestep2[20]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[4]~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[4]~28 .extended_lut = "off";
defparam \M_rot[4]~28 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[4]~28 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~28 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_mask[4]~q ),
	.datac(!\M_rot_pass1~q ),
	.datad(!\M_rot_sel_fill1~q ),
	.datae(!\M_rot[4]~28_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~28 .extended_lut = "off";
defparam \A_shift_rot_result~28 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~28 .shared_arith = "off";

dffeas \A_shift_rot_result[12] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~28_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_shift_rot_result[12]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[12] .is_wysiwyg = "true";
defparam \A_shift_rot_result[12] .power_up = "low";

dffeas \M_pc_plus_one[10] (
	.clk(clk_clk),
	.d(\Add7~45_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_pc_plus_one[10]~q ),
	.prn(vcc));
defparam \M_pc_plus_one[10] .is_wysiwyg = "true";
defparam \M_pc_plus_one[10] .power_up = "low";

dffeas \A_inst_result[12] (
	.clk(clk_clk),
	.d(\M_pc_plus_one[10]~q ),
	.asdata(\M_alu_result[12]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\A_inst_result[9]~0_combout ),
	.sload(!\M_exc_any~combout ),
	.ena(!\A_mem_stall~q ),
	.q(\A_inst_result[12]~q ),
	.prn(vcc));
defparam \A_inst_result[12] .is_wysiwyg = "true";
defparam \A_inst_result[12] .power_up = "low";

dffeas \A_mul_cell_p1[12] (
	.clk(clk_clk),
	.d(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[12]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_mul_cell_p1[12]~q ),
	.prn(vcc));
defparam \A_mul_cell_p1[12] .is_wysiwyg = "true";
defparam \A_mul_cell_p1[12] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[12]~30 (
	.dataa(!\A_slow_inst_result[12]~q ),
	.datab(!\A_shift_rot_result[12]~q ),
	.datac(!\A_inst_result[12]~q ),
	.datad(!\A_mul_cell_p1[12]~q ),
	.datae(!\A_wr_data_unfiltered[15]~0_combout ),
	.dataf(!\A_wr_data_unfiltered[15]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[12]~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[12]~30 .extended_lut = "off";
defparam \A_wr_data_unfiltered[12]~30 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_wr_data_unfiltered[12]~30 .shared_arith = "off";

dffeas \W_wr_data[12] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[12]~30_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[12]~q ),
	.prn(vcc));
defparam \W_wr_data[12] .is_wysiwyg = "true";
defparam \W_wr_data[12] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[12]~64 (
	.dataa(!\D_src2_reg[0]~7_combout ),
	.datab(!\D_src2_reg[0]~8_combout ),
	.datac(!\W_wr_data[12]~q ),
	.datad(!\A_wr_data_unfiltered[12]~30_combout ),
	.datae(!\M_alu_result[12]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[12]~64_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[12]~64 .extended_lut = "off";
defparam \D_src2_reg[12]~64 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \D_src2_reg[12]~64 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[12]~65 (
	.dataa(!\D_src2_reg[0]~4_combout ),
	.datab(!\D_src2_reg[0]~5_combout ),
	.datac(!\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[12] ),
	.datad(!\E_alu_result[12]~combout ),
	.datae(!\D_src2_reg[12]~64_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[12]~65_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[12]~65 .extended_lut = "off";
defparam \D_src2_reg[12]~65 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \D_src2_reg[12]~65 .shared_arith = "off";

dffeas \E_src2[12] (
	.clk(clk_clk),
	.d(\D_iw[18]~q ),
	.asdata(\D_src2_reg[12]~65_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src2[5]~2_combout ),
	.sload(!\D_ctrl_src2_choose_imm~q ),
	.ena(!\A_mem_stall~q ),
	.q(\E_src2[12]~q ),
	.prn(vcc));
defparam \E_src2[12] .is_wysiwyg = "true";
defparam \E_src2[12] .power_up = "low";

cyclonev_lcell_comb \E_alu_result~21 (
	.dataa(!\E_src2[12]~q ),
	.datab(!\E_src1[12]~q ),
	.datac(!\E_logic_op[1]~q ),
	.datad(!\E_logic_op[0]~q ),
	.datae(!\E_ctrl_logic~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result~21 .extended_lut = "off";
defparam \E_alu_result~21 .lut_mask = 64'h6996FFFF6996FFFF;
defparam \E_alu_result~21 .shared_arith = "off";

dffeas \E_extra_pc[10] (
	.clk(clk_clk),
	.d(\Add1~9_sumout ),
	.asdata(\D_pc_plus_one[10]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_br_pred_not_taken~combout ),
	.ena(!\A_mem_stall~q ),
	.q(\E_extra_pc[10]~q ),
	.prn(vcc));
defparam \E_extra_pc[10] .is_wysiwyg = "true";
defparam \E_extra_pc[10] .power_up = "low";

cyclonev_lcell_comb \E_alu_result[12] (
	.dataa(!\Add9~29_sumout ),
	.datab(!\E_ctrl_retaddr~q ),
	.datac(!\E_alu_result~0_combout ),
	.datad(!\E_alu_result~21_combout ),
	.datae(!\E_extra_pc[10]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[12]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[12] .extended_lut = "off";
defparam \E_alu_result[12] .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \E_alu_result[12] .shared_arith = "off";

dffeas \M_alu_result[12] (
	.clk(clk_clk),
	.d(\E_alu_result[12]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_alu_result[12]~q ),
	.prn(vcc));
defparam \M_alu_result[12] .is_wysiwyg = "true";
defparam \M_alu_result[12] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[12]~28 (
	.dataa(!\M_alu_result[12]~q ),
	.datab(!\A_wr_data_unfiltered[12]~30_combout ),
	.datac(!\first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[12] ),
	.datad(!\W_wr_data[12]~q ),
	.datae(!\E_src1[26]~0_combout ),
	.dataf(!\E_src1[26]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[12]~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[12]~28 .extended_lut = "off";
defparam \D_src1_reg[12]~28 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[12]~28 .shared_arith = "off";

dffeas \E_src1[12] (
	.clk(clk_clk),
	.d(\D_src1_reg[12]~28_combout ),
	.asdata(\E_alu_result[12]~combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\Equal303~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(!\A_mem_stall~q ),
	.q(\E_src1[12]~q ),
	.prn(vcc));
defparam \E_src1[12] .is_wysiwyg = "true";
defparam \E_src1[12] .power_up = "low";

cyclonev_lcell_comb \E_rot_step1[12]~4 (
	.dataa(!\E_src1[12]~q ),
	.datab(!\E_src1[11]~q ),
	.datac(!\E_src1[10]~q ),
	.datad(!\E_src1[9]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add10~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[12]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[12]~4 .extended_lut = "off";
defparam \E_rot_step1[12]~4 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[12]~4 .shared_arith = "off";

dffeas \M_rot_prestep2[16] (
	.clk(clk_clk),
	.d(\E_rot_step1[12]~4_combout ),
	.asdata(\E_rot_step1[16]~5_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add10~1_combout ),
	.ena(!\A_mem_stall~q ),
	.q(\M_rot_prestep2[16]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[16] .is_wysiwyg = "true";
defparam \M_rot_prestep2[16] .power_up = "low";

cyclonev_lcell_comb \M_rot[0]~26 (
	.dataa(!\M_rot_prestep2[16]~q ),
	.datab(!\M_rot_prestep2[8]~q ),
	.datac(!\M_rot_prestep2[0]~q ),
	.datad(!\M_rot_prestep2[24]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[0]~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[0]~26 .extended_lut = "off";
defparam \M_rot[0]~26 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[0]~26 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~26 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_mask[0]~q ),
	.datac(!\M_rot_pass2~q ),
	.datad(!\M_rot_sel_fill2~q ),
	.datae(!\M_rot[0]~26_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~26 .extended_lut = "off";
defparam \A_shift_rot_result~26 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~26 .shared_arith = "off";

dffeas \A_shift_rot_result[16] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~26_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_shift_rot_result[16]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[16] .is_wysiwyg = "true";
defparam \A_shift_rot_result[16] .power_up = "low";

dffeas \E_pc[14] (
	.clk(clk_clk),
	.d(\D_pc[14]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_pc[14]~q ),
	.prn(vcc));
defparam \E_pc[14] .is_wysiwyg = "true";
defparam \E_pc[14] .power_up = "low";

cyclonev_lcell_comb \Add7~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_pc[14]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add7~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add7~37_sumout ),
	.cout(),
	.shareout());
defparam \Add7~37 .extended_lut = "off";
defparam \Add7~37 .lut_mask = 64'h00000000000000FF;
defparam \Add7~37 .shared_arith = "off";

dffeas \M_pc_plus_one[14] (
	.clk(clk_clk),
	.d(\Add7~37_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_pc_plus_one[14]~q ),
	.prn(vcc));
defparam \M_pc_plus_one[14] .is_wysiwyg = "true";
defparam \M_pc_plus_one[14] .power_up = "low";

dffeas \E_iw[9] (
	.clk(clk_clk),
	.d(\D_iw[9]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_iw[9]~q ),
	.prn(vcc));
defparam \E_iw[9] .is_wysiwyg = "true";
defparam \E_iw[9] .power_up = "low";

dffeas \E_iw[7] (
	.clk(clk_clk),
	.d(\D_iw[7]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_iw[7]~q ),
	.prn(vcc));
defparam \E_iw[7] .is_wysiwyg = "true";
defparam \E_iw[7] .power_up = "low";

dffeas \E_iw[6] (
	.clk(clk_clk),
	.d(\D_iw[6]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_iw[6]~q ),
	.prn(vcc));
defparam \E_iw[6] .is_wysiwyg = "true";
defparam \E_iw[6] .power_up = "low";

dffeas \E_iw[10] (
	.clk(clk_clk),
	.d(\D_iw[10]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_iw[10]~q ),
	.prn(vcc));
defparam \E_iw[10] .is_wysiwyg = "true";
defparam \E_iw[10] .power_up = "low";

dffeas \E_iw[8] (
	.clk(clk_clk),
	.d(\D_iw[8]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_iw[8]~q ),
	.prn(vcc));
defparam \E_iw[8] .is_wysiwyg = "true";
defparam \E_iw[8] .power_up = "low";

cyclonev_lcell_comb \M_control_reg_rddata[16]~0 (
	.dataa(!\E_iw[9]~q ),
	.datab(!\E_iw[7]~q ),
	.datac(!\E_iw[6]~q ),
	.datad(!\E_iw[10]~q ),
	.datae(!\E_iw[8]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_control_reg_rddata[16]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_control_reg_rddata[16]~0 .extended_lut = "off";
defparam \M_control_reg_rddata[16]~0 .lut_mask = 64'hFF96FFFFFF96FFFF;
defparam \M_control_reg_rddata[16]~0 .shared_arith = "off";

dffeas \M_iw[7] (
	.clk(clk_clk),
	.d(\E_iw[7]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_iw[7]~q ),
	.prn(vcc));
defparam \M_iw[7] .is_wysiwyg = "true";
defparam \M_iw[7] .power_up = "low";

dffeas \A_iw[7] (
	.clk(clk_clk),
	.d(\M_iw[7]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_iw[7]~q ),
	.prn(vcc));
defparam \A_iw[7] .is_wysiwyg = "true";
defparam \A_iw[7] .power_up = "low";

dffeas \M_iw[6] (
	.clk(clk_clk),
	.d(\E_iw[6]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_iw[6]~q ),
	.prn(vcc));
defparam \M_iw[6] .is_wysiwyg = "true";
defparam \M_iw[6] .power_up = "low";

dffeas \A_iw[6] (
	.clk(clk_clk),
	.d(\M_iw[6]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_iw[6]~q ),
	.prn(vcc));
defparam \A_iw[6] .is_wysiwyg = "true";
defparam \A_iw[6] .power_up = "low";

dffeas \M_iw[10] (
	.clk(clk_clk),
	.d(\E_iw[10]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_iw[10]~q ),
	.prn(vcc));
defparam \M_iw[10] .is_wysiwyg = "true";
defparam \M_iw[10] .power_up = "low";

dffeas \A_iw[10] (
	.clk(clk_clk),
	.d(\M_iw[10]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_iw[10]~q ),
	.prn(vcc));
defparam \A_iw[10] .is_wysiwyg = "true";
defparam \A_iw[10] .power_up = "low";

dffeas \M_iw[9] (
	.clk(clk_clk),
	.d(\E_iw[9]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_iw[9]~q ),
	.prn(vcc));
defparam \M_iw[9] .is_wysiwyg = "true";
defparam \M_iw[9] .power_up = "low";

dffeas \A_iw[9] (
	.clk(clk_clk),
	.d(\M_iw[9]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_iw[9]~q ),
	.prn(vcc));
defparam \A_iw[9] .is_wysiwyg = "true";
defparam \A_iw[9] .power_up = "low";

dffeas \M_iw[8] (
	.clk(clk_clk),
	.d(\E_iw[8]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_iw[8]~q ),
	.prn(vcc));
defparam \M_iw[8] .is_wysiwyg = "true";
defparam \M_iw[8] .power_up = "low";

dffeas \A_iw[8] (
	.clk(clk_clk),
	.d(\M_iw[8]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_iw[8]~q ),
	.prn(vcc));
defparam \A_iw[8] .is_wysiwyg = "true";
defparam \A_iw[8] .power_up = "low";

cyclonev_lcell_comb E_op_wrctl(
	.dataa(!\E_iw[14]~q ),
	.datab(!\E_op_rdctl~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_op_wrctl~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam E_op_wrctl.extended_lut = "off";
defparam E_op_wrctl.lut_mask = 64'h7777777777777777;
defparam E_op_wrctl.shared_arith = "off";

dffeas M_ctrl_wrctl_inst(
	.clk(clk_clk),
	.d(\E_op_wrctl~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_ctrl_wrctl_inst~q ),
	.prn(vcc));
defparam M_ctrl_wrctl_inst.is_wysiwyg = "true";
defparam M_ctrl_wrctl_inst.power_up = "low";

dffeas A_ctrl_wrctl_inst(
	.clk(clk_clk),
	.d(\M_ctrl_wrctl_inst~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_ctrl_wrctl_inst~q ),
	.prn(vcc));
defparam A_ctrl_wrctl_inst.is_wysiwyg = "true";
defparam A_ctrl_wrctl_inst.power_up = "low";

cyclonev_lcell_comb \A_wrctl_status~0 (
	.dataa(!\A_iw[10]~q ),
	.datab(!\A_iw[9]~q ),
	.datac(!\A_iw[8]~q ),
	.datad(!\A_ctrl_wrctl_inst~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wrctl_status~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wrctl_status~0 .extended_lut = "off";
defparam \A_wrctl_status~0 .lut_mask = 64'hFEFFFEFFFEFFFEFF;
defparam \A_wrctl_status~0 .shared_arith = "off";

cyclonev_lcell_comb \W_ienable_reg_irq1_nxt~0 (
	.dataa(!\A_valid_from_M~q ),
	.datab(!\A_iw[7]~q ),
	.datac(!\A_iw[6]~q ),
	.datad(!\A_wrctl_status~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_ienable_reg_irq1_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_ienable_reg_irq1_nxt~0 .extended_lut = "off";
defparam \W_ienable_reg_irq1_nxt~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \W_ienable_reg_irq1_nxt~0 .shared_arith = "off";

dffeas W_ienable_reg_irq16(
	.clk(clk_clk),
	.d(\A_inst_result[16]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_ienable_reg_irq1_nxt~0_combout ),
	.q(\W_ienable_reg_irq16~q ),
	.prn(vcc));
defparam W_ienable_reg_irq16.is_wysiwyg = "true";
defparam W_ienable_reg_irq16.power_up = "low";

cyclonev_lcell_comb \W_ipending_reg_irq16_nxt~0 (
	.dataa(!\W_ienable_reg_irq16~q ),
	.datab(!\the_first_nios2_system_cpu_cpu_nios2_oci|the_first_nios2_system_cpu_cpu_nios2_avalon_reg|oci_ienable[16]~q ),
	.datac(!av_readdata_9),
	.datad(!av_readdata_8),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_ipending_reg_irq16_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_ipending_reg_irq16_nxt~0 .extended_lut = "off";
defparam \W_ipending_reg_irq16_nxt~0 .lut_mask = 64'hDFFFDFFFDFFFDFFF;
defparam \W_ipending_reg_irq16_nxt~0 .shared_arith = "off";

dffeas W_ipending_reg_irq16(
	.clk(clk_clk),
	.d(\W_ipending_reg_irq16_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_ipending_reg_irq16~q ),
	.prn(vcc));
defparam W_ipending_reg_irq16.is_wysiwyg = "true";
defparam W_ipending_reg_irq16.power_up = "low";

cyclonev_lcell_comb \Equal324~0 (
	.dataa(!\D_iw[10]~q ),
	.datab(!\D_iw[6]~q ),
	.datac(!\D_iw[7]~q ),
	.datad(!\D_iw[8]~q ),
	.datae(!\D_iw[9]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal324~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal324~0 .extended_lut = "off";
defparam \Equal324~0 .lut_mask = 64'hFFFFFFBFFFFFFFBF;
defparam \Equal324~0 .shared_arith = "off";

cyclonev_lcell_comb \E_control_reg_rddata[1]~0 (
	.dataa(!\D_iw[10]~q ),
	.datab(!\D_iw[6]~q ),
	.datac(!\D_iw[7]~q ),
	.datad(!\D_iw[8]~q ),
	.datae(!\D_iw[9]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_control_reg_rddata[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_control_reg_rddata[1]~0 .extended_lut = "off";
defparam \E_control_reg_rddata[1]~0 .lut_mask = 64'hFFFFEBBEFFFFEBBE;
defparam \E_control_reg_rddata[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \D_control_reg_rddata_muxed[16]~3 (
	.dataa(!\W_ipending_reg_irq16~q ),
	.datab(!\W_ienable_reg_irq16~q ),
	.datac(!\Equal324~0_combout ),
	.datad(!\E_control_reg_rddata[1]~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_control_reg_rddata_muxed[16]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_control_reg_rddata_muxed[16]~3 .extended_lut = "off";
defparam \D_control_reg_rddata_muxed[16]~3 .lut_mask = 64'h53FF53FF53FF53FF;
defparam \D_control_reg_rddata_muxed[16]~3 .shared_arith = "off";

dffeas \E_control_reg_rddata[16] (
	.clk(clk_clk),
	.d(\D_control_reg_rddata_muxed[16]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_control_reg_rddata[16]~q ),
	.prn(vcc));
defparam \E_control_reg_rddata[16] .is_wysiwyg = "true";
defparam \E_control_reg_rddata[16] .power_up = "low";

cyclonev_lcell_comb \E_control_reg_rddata_muxed[16]~5 (
	.dataa(!\M_control_reg_rddata[16]~0_combout ),
	.datab(!\E_control_reg_rddata[16]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_control_reg_rddata_muxed[16]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_control_reg_rddata_muxed[16]~5 .extended_lut = "off";
defparam \E_control_reg_rddata_muxed[16]~5 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \E_control_reg_rddata_muxed[16]~5 .shared_arith = "off";

dffeas \M_control_reg_rddata[16] (
	.clk(clk_clk),
	.d(\E_control_reg_rddata_muxed[16]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_control_reg_rddata[16]~q ),
	.prn(vcc));
defparam \M_control_reg_rddata[16] .is_wysiwyg = "true";
defparam \M_control_reg_rddata[16] .power_up = "low";

cyclonev_lcell_comb \M_inst_result[16]~5 (
	.dataa(!\M_exc_any~combout ),
	.datab(!\M_alu_result[16]~q ),
	.datac(!\M_ctrl_rd_ctl_reg~q ),
	.datad(!\M_pc_plus_one[14]~q ),
	.datae(!\M_control_reg_rddata[16]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_inst_result[16]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_inst_result[16]~5 .extended_lut = "off";
defparam \M_inst_result[16]~5 .lut_mask = 64'h7BFFFFFF7BFFFFFF;
defparam \M_inst_result[16]~5 .shared_arith = "off";

dffeas \A_inst_result[16] (
	.clk(clk_clk),
	.d(\M_inst_result[16]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_inst_result[16]~q ),
	.prn(vcc));
defparam \A_inst_result[16] .is_wysiwyg = "true";
defparam \A_inst_result[16] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[16]~28 (
	.dataa(!\A_slow_inst_result[16]~q ),
	.datab(!\A_shift_rot_result[16]~q ),
	.datac(!\A_inst_result[16]~q ),
	.datad(!\Add12~57_sumout ),
	.datae(!\A_wr_data_unfiltered[15]~0_combout ),
	.dataf(!\A_wr_data_unfiltered[15]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[16]~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[16]~28 .extended_lut = "off";
defparam \A_wr_data_unfiltered[16]~28 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_wr_data_unfiltered[16]~28 .shared_arith = "off";

dffeas \W_wr_data[16] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[16]~28_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[16]~q ),
	.prn(vcc));
defparam \W_wr_data[16] .is_wysiwyg = "true";
defparam \W_wr_data[16] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[16]~61 (
	.dataa(!\D_src2_reg[0]~4_combout ),
	.datab(!\D_src2_reg[0]~7_combout ),
	.datac(!\D_src2_reg[0]~8_combout ),
	.datad(!\M_alu_result[16]~q ),
	.datae(!\A_wr_data_unfiltered[16]~28_combout ),
	.dataf(!\W_wr_data[16]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[16]~61_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[16]~61 .extended_lut = "off";
defparam \D_src2_reg[16]~61 .lut_mask = 64'hBEFFFFFFFFFFFFFF;
defparam \D_src2_reg[16]~61 .shared_arith = "off";

cyclonev_lcell_comb \E_logic_result[16]~12 (
	.dataa(!\E_src2[16]~q ),
	.datab(!\E_src1[16]~q ),
	.datac(!\E_logic_op[1]~q ),
	.datad(!\E_logic_op[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[16]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[16]~12 .extended_lut = "off";
defparam \E_logic_result[16]~12 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[16]~12 .shared_arith = "off";

dffeas \E_extra_pc[14] (
	.clk(clk_clk),
	.d(\Add1~1_sumout ),
	.asdata(\D_pc_plus_one[14]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_br_pred_not_taken~combout ),
	.ena(!\A_mem_stall~q ),
	.q(\E_extra_pc[14]~q ),
	.prn(vcc));
defparam \E_extra_pc[14] .is_wysiwyg = "true";
defparam \E_extra_pc[14] .power_up = "low";

cyclonev_lcell_comb \E_alu_result[16]~19 (
	.dataa(!\E_logic_result[16]~12_combout ),
	.datab(!\E_ctrl_logic~q ),
	.datac(!\E_ctrl_retaddr~q ),
	.datad(!\E_extra_pc[14]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[16]~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[16]~19 .extended_lut = "off";
defparam \E_alu_result[16]~19 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \E_alu_result[16]~19 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[16]~31 (
	.dataa(!\D_ctrl_hi_imm16~q ),
	.datab(!\D_iw[21]~q ),
	.datac(!\D_ctrl_unsigned_lo_imm16~q ),
	.datad(!\D_iw[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[16]~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[16]~31 .extended_lut = "off";
defparam \D_src2[16]~31 .lut_mask = 64'h7BFF7BFF7BFF7BFF;
defparam \D_src2[16]~31 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[16]~32 (
	.dataa(!\D_ctrl_src2_choose_imm~q ),
	.datab(!\Add9~13_sumout ),
	.datac(!\E_alu_result~0_combout ),
	.datad(!\E_alu_result[16]~19_combout ),
	.datae(!\D_src2[16]~31_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[16]~32_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[16]~32 .extended_lut = "off";
defparam \D_src2[16]~32 .lut_mask = 64'hFFFFFFD8FFFFFFD8;
defparam \D_src2[16]~32 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[16]~26 (
	.dataa(!\D_src2_reg[0]~5_combout ),
	.datab(!\D_ctrl_src2_choose_imm~q ),
	.datac(!\D_src2_reg[16]~61_combout ),
	.datad(!\D_src2_reg[0]~4_combout ),
	.datae(!\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[16] ),
	.dataf(!\D_src2[16]~32_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[16]~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[16]~26 .extended_lut = "off";
defparam \D_src2[16]~26 .lut_mask = 64'hFFFFFFFF6FFFFFFF;
defparam \D_src2[16]~26 .shared_arith = "off";

dffeas \E_src2[16] (
	.clk(clk_clk),
	.d(\D_src2[16]~26_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src2[30]~1_combout ),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_src2[16]~q ),
	.prn(vcc));
defparam \E_src2[16] .is_wysiwyg = "true";
defparam \E_src2[16] .power_up = "low";

cyclonev_lcell_comb \E_alu_result[16] (
	.dataa(!\Add9~13_sumout ),
	.datab(!\E_alu_result~0_combout ),
	.datac(!\E_alu_result[16]~19_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[16]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[16] .extended_lut = "off";
defparam \E_alu_result[16] .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \E_alu_result[16] .shared_arith = "off";

dffeas \M_alu_result[16] (
	.clk(clk_clk),
	.d(\E_alu_result[16]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_alu_result[16]~q ),
	.prn(vcc));
defparam \M_alu_result[16] .is_wysiwyg = "true";
defparam \M_alu_result[16] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[16]~26 (
	.dataa(!\M_alu_result[16]~q ),
	.datab(!\A_wr_data_unfiltered[16]~28_combout ),
	.datac(!\first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[16] ),
	.datad(!\W_wr_data[16]~q ),
	.datae(!\E_src1[26]~0_combout ),
	.dataf(!\E_src1[26]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[16]~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[16]~26 .extended_lut = "off";
defparam \D_src1_reg[16]~26 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[16]~26 .shared_arith = "off";

dffeas \E_src1[16] (
	.clk(clk_clk),
	.d(\D_src1_reg[16]~26_combout ),
	.asdata(\E_alu_result[16]~combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\Equal303~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(!\A_mem_stall~q ),
	.q(\E_src1[16]~q ),
	.prn(vcc));
defparam \E_src1[16] .is_wysiwyg = "true";
defparam \E_src1[16] .power_up = "low";

cyclonev_lcell_comb \E_rot_step1[16]~5 (
	.dataa(!\E_src1[16]~q ),
	.datab(!\E_src1[15]~q ),
	.datac(!\E_src1[14]~q ),
	.datad(!\E_src1[13]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add10~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[16]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[16]~5 .extended_lut = "off";
defparam \E_rot_step1[16]~5 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[16]~5 .shared_arith = "off";

dffeas \M_rot_prestep2[20] (
	.clk(clk_clk),
	.d(\E_rot_step1[16]~5_combout ),
	.asdata(\E_rot_step1[20]~2_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add10~1_combout ),
	.ena(!\A_mem_stall~q ),
	.q(\M_rot_prestep2[20]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[20] .is_wysiwyg = "true";
defparam \M_rot_prestep2[20] .power_up = "low";

cyclonev_lcell_comb \M_rot[4]~21 (
	.dataa(!\M_rot_prestep2[20]~q ),
	.datab(!\M_rot_prestep2[12]~q ),
	.datac(!\M_rot_prestep2[4]~q ),
	.datad(!\M_rot_prestep2[28]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[4]~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[4]~21 .extended_lut = "off";
defparam \M_rot[4]~21 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[4]~21 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~21 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_mask[4]~q ),
	.datac(!\M_rot_pass2~q ),
	.datad(!\M_rot_sel_fill2~q ),
	.datae(!\M_rot[4]~21_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~21 .extended_lut = "off";
defparam \A_shift_rot_result~21 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~21 .shared_arith = "off";

dffeas \A_shift_rot_result[20] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~21_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_shift_rot_result[20]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[20] .is_wysiwyg = "true";
defparam \A_shift_rot_result[20] .power_up = "low";

dffeas \A_inst_result[20] (
	.clk(clk_clk),
	.d(\M_alu_result[20]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\A_inst_result[26]~1_combout ),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_inst_result[20]~q ),
	.prn(vcc));
defparam \A_inst_result[20] .is_wysiwyg = "true";
defparam \A_inst_result[20] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[20]~23 (
	.dataa(!\A_slow_inst_result[20]~q ),
	.datab(!\A_shift_rot_result[20]~q ),
	.datac(!\A_inst_result[20]~q ),
	.datad(!\Add12~37_sumout ),
	.datae(!\A_wr_data_unfiltered[15]~0_combout ),
	.dataf(!\A_wr_data_unfiltered[15]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[20]~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[20]~23 .extended_lut = "off";
defparam \A_wr_data_unfiltered[20]~23 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_wr_data_unfiltered[20]~23 .shared_arith = "off";

dffeas \W_wr_data[20] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[20]~23_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[20]~q ),
	.prn(vcc));
defparam \W_wr_data[20] .is_wysiwyg = "true";
defparam \W_wr_data[20] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[20]~54 (
	.dataa(!\D_src2_reg[0]~4_combout ),
	.datab(!\D_src2_reg[0]~7_combout ),
	.datac(!\D_src2_reg[0]~8_combout ),
	.datad(!\M_alu_result[20]~q ),
	.datae(!\A_wr_data_unfiltered[20]~23_combout ),
	.dataf(!\W_wr_data[20]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[20]~54_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[20]~54 .extended_lut = "off";
defparam \D_src2_reg[20]~54 .lut_mask = 64'hBEFFFFFFFFFFFFFF;
defparam \D_src2_reg[20]~54 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[20]~39 (
	.dataa(!\D_ctrl_hi_imm16~q ),
	.datab(!\D_iw[10]~q ),
	.datac(!\D_iw[21]~q ),
	.datad(!\D_ctrl_unsigned_lo_imm16~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[20]~39_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[20]~39 .extended_lut = "off";
defparam \D_src2[20]~39 .lut_mask = 64'h7FBF7FBF7FBF7FBF;
defparam \D_src2[20]~39 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[20]~40 (
	.dataa(!\D_ctrl_src2_choose_imm~q ),
	.datab(!\E_logic_result[20]~9_combout ),
	.datac(!\E_ctrl_logic~q ),
	.datad(!\E_alu_result~0_combout ),
	.datae(!\Add9~109_sumout ),
	.dataf(!\D_src2[20]~39_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[20]~40_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[20]~40 .extended_lut = "off";
defparam \D_src2[20]~40 .lut_mask = 64'h27FFFFFFFFFFFFFF;
defparam \D_src2[20]~40 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[20]~19 (
	.dataa(!\D_src2_reg[0]~5_combout ),
	.datab(!\D_ctrl_src2_choose_imm~q ),
	.datac(!\D_src2_reg[20]~54_combout ),
	.datad(!\D_src2_reg[0]~4_combout ),
	.datae(!\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[20] ),
	.dataf(!\D_src2[20]~40_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[20]~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[20]~19 .extended_lut = "off";
defparam \D_src2[20]~19 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \D_src2[20]~19 .shared_arith = "off";

dffeas \E_src2[20] (
	.clk(clk_clk),
	.d(\D_src2[20]~19_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src2[30]~1_combout ),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_src2[20]~q ),
	.prn(vcc));
defparam \E_src2[20] .is_wysiwyg = "true";
defparam \E_src2[20] .power_up = "low";

cyclonev_lcell_comb \E_logic_result[20]~9 (
	.dataa(!\E_src2[20]~q ),
	.datab(!\E_src1[20]~q ),
	.datac(!\E_logic_op[1]~q ),
	.datad(!\E_logic_op[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[20]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[20]~9 .extended_lut = "off";
defparam \E_logic_result[20]~9 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[20]~9 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[20] (
	.dataa(!\E_logic_result[20]~9_combout ),
	.datab(!\E_ctrl_logic~q ),
	.datac(!\E_alu_result~0_combout ),
	.datad(!\Add9~109_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[20]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[20] .extended_lut = "off";
defparam \E_alu_result[20] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \E_alu_result[20] .shared_arith = "off";

dffeas \M_alu_result[20] (
	.clk(clk_clk),
	.d(\E_alu_result[20]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_alu_result[20]~q ),
	.prn(vcc));
defparam \M_alu_result[20] .is_wysiwyg = "true";
defparam \M_alu_result[20] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[20]~20 (
	.dataa(!\M_alu_result[20]~q ),
	.datab(!\A_wr_data_unfiltered[20]~23_combout ),
	.datac(!\first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[20] ),
	.datad(!\W_wr_data[20]~q ),
	.datae(!\E_src1[26]~0_combout ),
	.dataf(!\E_src1[26]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[20]~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[20]~20 .extended_lut = "off";
defparam \D_src1_reg[20]~20 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[20]~20 .shared_arith = "off";

dffeas \E_src1[20] (
	.clk(clk_clk),
	.d(\D_src1_reg[20]~20_combout ),
	.asdata(\E_alu_result[20]~combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\Equal303~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(!\A_mem_stall~q ),
	.q(\E_src1[20]~q ),
	.prn(vcc));
defparam \E_src1[20] .is_wysiwyg = "true";
defparam \E_src1[20] .power_up = "low";

cyclonev_lcell_comb \E_rot_step1[20]~2 (
	.dataa(!\E_src1[20]~q ),
	.datab(!\E_src1[19]~q ),
	.datac(!\E_src1[18]~q ),
	.datad(!\E_src1[17]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add10~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[20]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[20]~2 .extended_lut = "off";
defparam \E_rot_step1[20]~2 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[20]~2 .shared_arith = "off";

dffeas \M_rot_prestep2[24] (
	.clk(clk_clk),
	.d(\E_rot_step1[20]~2_combout ),
	.asdata(\E_rot_step1[24]~3_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add10~1_combout ),
	.ena(!\A_mem_stall~q ),
	.q(\M_rot_prestep2[24]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[24] .is_wysiwyg = "true";
defparam \M_rot_prestep2[24] .power_up = "low";

cyclonev_lcell_comb \M_rot[0]~18 (
	.dataa(!\M_rot_prestep2[8]~q ),
	.datab(!\M_rot_prestep2[0]~q ),
	.datac(!\M_rot_prestep2[24]~q ),
	.datad(!\M_rot_prestep2[16]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[0]~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[0]~18 .extended_lut = "off";
defparam \M_rot[0]~18 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[0]~18 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~18 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_mask[0]~q ),
	.datac(!\M_rot_pass1~q ),
	.datad(!\M_rot_sel_fill1~q ),
	.datae(!\M_rot[0]~18_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~18 .extended_lut = "off";
defparam \A_shift_rot_result~18 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~18 .shared_arith = "off";

dffeas \A_shift_rot_result[8] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~18_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_shift_rot_result[8]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[8] .is_wysiwyg = "true";
defparam \A_shift_rot_result[8] .power_up = "low";

dffeas \M_pc_plus_one[6] (
	.clk(clk_clk),
	.d(\Add7~29_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_pc_plus_one[6]~q ),
	.prn(vcc));
defparam \M_pc_plus_one[6] .is_wysiwyg = "true";
defparam \M_pc_plus_one[6] .power_up = "low";

dffeas \A_inst_result[8] (
	.clk(clk_clk),
	.d(\M_pc_plus_one[6]~q ),
	.asdata(\M_alu_result[8]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\A_inst_result[9]~0_combout ),
	.sload(!\M_exc_any~combout ),
	.ena(!\A_mem_stall~q ),
	.q(\A_inst_result[8]~q ),
	.prn(vcc));
defparam \A_inst_result[8] .is_wysiwyg = "true";
defparam \A_inst_result[8] .power_up = "low";

dffeas \A_mul_cell_p1[8] (
	.clk(clk_clk),
	.d(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[8]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_mul_cell_p1[8]~q ),
	.prn(vcc));
defparam \A_mul_cell_p1[8] .is_wysiwyg = "true";
defparam \A_mul_cell_p1[8] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[8]~20 (
	.dataa(!\A_slow_inst_result[8]~q ),
	.datab(!\A_shift_rot_result[8]~q ),
	.datac(!\A_inst_result[8]~q ),
	.datad(!\A_mul_cell_p1[8]~q ),
	.datae(!\A_wr_data_unfiltered[15]~0_combout ),
	.dataf(!\A_wr_data_unfiltered[15]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[8]~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[8]~20 .extended_lut = "off";
defparam \A_wr_data_unfiltered[8]~20 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_wr_data_unfiltered[8]~20 .shared_arith = "off";

dffeas \W_wr_data[8] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[8]~20_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[8]~q ),
	.prn(vcc));
defparam \W_wr_data[8] .is_wysiwyg = "true";
defparam \W_wr_data[8] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[8]~48 (
	.dataa(!\D_src2_reg[0]~7_combout ),
	.datab(!\D_src2_reg[0]~8_combout ),
	.datac(!\W_wr_data[8]~q ),
	.datad(!\A_wr_data_unfiltered[8]~20_combout ),
	.datae(!\M_alu_result[8]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[8]~48_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[8]~48 .extended_lut = "off";
defparam \D_src2_reg[8]~48 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \D_src2_reg[8]~48 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[8]~49 (
	.dataa(!\D_src2_reg[0]~4_combout ),
	.datab(!\D_src2_reg[0]~5_combout ),
	.datac(!\D_src2_reg[8]~48_combout ),
	.datad(!\E_alu_result[8]~combout ),
	.datae(!\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[8] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[8]~49_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[8]~49 .extended_lut = "off";
defparam \D_src2_reg[8]~49 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \D_src2_reg[8]~49 .shared_arith = "off";

dffeas \E_src2[8] (
	.clk(clk_clk),
	.d(\D_iw[14]~q ),
	.asdata(\D_src2_reg[8]~49_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src2[5]~2_combout ),
	.sload(!\D_ctrl_src2_choose_imm~q ),
	.ena(!\A_mem_stall~q ),
	.q(\E_src2[8]~q ),
	.prn(vcc));
defparam \E_src2[8] .is_wysiwyg = "true";
defparam \E_src2[8] .power_up = "low";

cyclonev_lcell_comb \E_alu_result~15 (
	.dataa(!\E_src2[8]~q ),
	.datab(!\E_src1[8]~q ),
	.datac(!\E_logic_op[1]~q ),
	.datad(!\E_logic_op[0]~q ),
	.datae(!\E_ctrl_logic~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result~15 .extended_lut = "off";
defparam \E_alu_result~15 .lut_mask = 64'h6996FFFF6996FFFF;
defparam \E_alu_result~15 .shared_arith = "off";

dffeas \D_pc_plus_one[6] (
	.clk(clk_clk),
	.d(\Add3~25_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_pc_plus_one[6]~q ),
	.prn(vcc));
defparam \D_pc_plus_one[6] .is_wysiwyg = "true";
defparam \D_pc_plus_one[6] .power_up = "low";

dffeas \E_extra_pc[6] (
	.clk(clk_clk),
	.d(\D_br_taken_waddr_partial[6]~q ),
	.asdata(\D_pc_plus_one[6]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_br_pred_not_taken~combout ),
	.ena(!\A_mem_stall~q ),
	.q(\E_extra_pc[6]~q ),
	.prn(vcc));
defparam \E_extra_pc[6] .is_wysiwyg = "true";
defparam \E_extra_pc[6] .power_up = "low";

cyclonev_lcell_comb \E_alu_result[8] (
	.dataa(!\Add9~9_sumout ),
	.datab(!\E_ctrl_retaddr~q ),
	.datac(!\E_alu_result~0_combout ),
	.datad(!\E_alu_result~15_combout ),
	.datae(!\E_extra_pc[6]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[8]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[8] .extended_lut = "off";
defparam \E_alu_result[8] .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \E_alu_result[8] .shared_arith = "off";

dffeas \M_alu_result[8] (
	.clk(clk_clk),
	.d(\E_alu_result[8]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_alu_result[8]~q ),
	.prn(vcc));
defparam \M_alu_result[8] .is_wysiwyg = "true";
defparam \M_alu_result[8] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[8]~14 (
	.dataa(!\M_alu_result[8]~q ),
	.datab(!\A_wr_data_unfiltered[8]~20_combout ),
	.datac(!\first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[8] ),
	.datad(!\W_wr_data[8]~q ),
	.datae(!\E_src1[26]~0_combout ),
	.dataf(!\E_src1[26]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[8]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[8]~14 .extended_lut = "off";
defparam \D_src1_reg[8]~14 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[8]~14 .shared_arith = "off";

dffeas \E_src1[8] (
	.clk(clk_clk),
	.d(\D_src1_reg[8]~14_combout ),
	.asdata(\E_alu_result[8]~combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\Equal303~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(!\A_mem_stall~q ),
	.q(\E_src1[8]~q ),
	.prn(vcc));
defparam \E_src1[8] .is_wysiwyg = "true";
defparam \E_src1[8] .power_up = "low";

dffeas \M_target_pcb[8] (
	.clk(clk_clk),
	.d(\E_src1[8]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_target_pcb[8]~q ),
	.prn(vcc));
defparam \M_target_pcb[8] .is_wysiwyg = "true";
defparam \M_target_pcb[8] .power_up = "low";

cyclonev_lcell_comb \A_pipe_flush_waddr_nxt~6 (
	.dataa(!\M_exc_any~combout ),
	.datab(!\M_pc_plus_one[6]~q ),
	.datac(!\M_ctrl_jmp_indirect~q ),
	.datad(!\M_target_pcb[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_pipe_flush_waddr_nxt~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_pipe_flush_waddr_nxt~6 .extended_lut = "off";
defparam \A_pipe_flush_waddr_nxt~6 .lut_mask = 64'hA3FFA3FFA3FFA3FF;
defparam \A_pipe_flush_waddr_nxt~6 .shared_arith = "off";

dffeas \A_pipe_flush_waddr[6] (
	.clk(clk_clk),
	.d(\A_pipe_flush_waddr_nxt~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\M_exc_break~0_combout ),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_pipe_flush_waddr[6]~q ),
	.prn(vcc));
defparam \A_pipe_flush_waddr[6] .is_wysiwyg = "true";
defparam \A_pipe_flush_waddr[6] .power_up = "low";

dffeas \M_pipe_flush_waddr[6] (
	.clk(clk_clk),
	.d(\E_extra_pc[6]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_pipe_flush_waddr[6]~q ),
	.prn(vcc));
defparam \M_pipe_flush_waddr[6] .is_wysiwyg = "true";
defparam \M_pipe_flush_waddr[6] .power_up = "low";

cyclonev_lcell_comb \F_ic_tag_rd_addr_nxt[3]~11 (
	.dataa(!\F_ic_tag_rd_addr_nxt[3]~10_combout ),
	.datab(!\E_src1[8]~q ),
	.datac(!\A_pipe_flush_waddr[6]~q ),
	.datad(!\M_pipe_flush_waddr[6]~q ),
	.datae(!\F_ic_tag_rd_addr_nxt[3]~2_combout ),
	.dataf(!\F_ic_tag_rd_addr_nxt[3]~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_tag_rd_addr_nxt[3]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_tag_rd_addr_nxt[3]~11 .extended_lut = "off";
defparam \F_ic_tag_rd_addr_nxt[3]~11 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \F_ic_tag_rd_addr_nxt[3]~11 .shared_arith = "off";

dffeas \F_pc[6] (
	.clk(clk_clk),
	.d(\F_ic_tag_rd_addr_nxt[3]~11_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\F_pc[6]~q ),
	.prn(vcc));
defparam \F_pc[6] .is_wysiwyg = "true";
defparam \F_pc[6] .power_up = "low";

cyclonev_lcell_comb \Add3~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\F_pc[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~29_sumout ),
	.cout(\Add3~30 ),
	.shareout());
defparam \Add3~29 .extended_lut = "off";
defparam \Add3~29 .lut_mask = 64'h00000000000000FF;
defparam \Add3~29 .shared_arith = "off";

cyclonev_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[15] ),
	.datae(gnd),
	.dataf(!\Add3~29_sumout ),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout());
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~37 .shared_arith = "off";

dffeas \D_br_taken_waddr_partial[7] (
	.clk(clk_clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_br_taken_waddr_partial[7]~q ),
	.prn(vcc));
defparam \D_br_taken_waddr_partial[7] .is_wysiwyg = "true";
defparam \D_br_taken_waddr_partial[7] .power_up = "low";

cyclonev_lcell_comb \F_ic_tag_rd_addr_nxt[4]~12 (
	.dataa(!\D_pc[7]~q ),
	.datab(!\D_br_taken_waddr_partial[7]~q ),
	.datac(!\Add3~29_sumout ),
	.datad(!\D_iw[13]~q ),
	.datae(!\F_ic_tag_rd_addr_nxt[3]~0_combout ),
	.dataf(!\F_ic_tag_rd_addr_nxt[3]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_tag_rd_addr_nxt[4]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_tag_rd_addr_nxt[4]~12 .extended_lut = "off";
defparam \F_ic_tag_rd_addr_nxt[4]~12 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \F_ic_tag_rd_addr_nxt[4]~12 .shared_arith = "off";

dffeas \M_target_pcb[9] (
	.clk(clk_clk),
	.d(\E_src1[9]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_target_pcb[9]~q ),
	.prn(vcc));
defparam \M_target_pcb[9] .is_wysiwyg = "true";
defparam \M_target_pcb[9] .power_up = "low";

cyclonev_lcell_comb \A_pipe_flush_waddr_nxt~7 (
	.dataa(!\M_exc_any~combout ),
	.datab(!\M_pc_plus_one[7]~q ),
	.datac(!\M_ctrl_jmp_indirect~q ),
	.datad(!\M_target_pcb[9]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_pipe_flush_waddr_nxt~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_pipe_flush_waddr_nxt~7 .extended_lut = "off";
defparam \A_pipe_flush_waddr_nxt~7 .lut_mask = 64'hA3FFA3FFA3FFA3FF;
defparam \A_pipe_flush_waddr_nxt~7 .shared_arith = "off";

dffeas \A_pipe_flush_waddr[7] (
	.clk(clk_clk),
	.d(\A_pipe_flush_waddr_nxt~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\M_exc_break~0_combout ),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_pipe_flush_waddr[7]~q ),
	.prn(vcc));
defparam \A_pipe_flush_waddr[7] .is_wysiwyg = "true";
defparam \A_pipe_flush_waddr[7] .power_up = "low";

dffeas \M_pipe_flush_waddr[7] (
	.clk(clk_clk),
	.d(\E_extra_pc[7]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_pipe_flush_waddr[7]~q ),
	.prn(vcc));
defparam \M_pipe_flush_waddr[7] .is_wysiwyg = "true";
defparam \M_pipe_flush_waddr[7] .power_up = "low";

cyclonev_lcell_comb \F_ic_tag_rd_addr_nxt[4]~13 (
	.dataa(!\F_ic_tag_rd_addr_nxt[4]~12_combout ),
	.datab(!\E_src1[9]~q ),
	.datac(!\A_pipe_flush_waddr[7]~q ),
	.datad(!\M_pipe_flush_waddr[7]~q ),
	.datae(!\F_ic_tag_rd_addr_nxt[3]~2_combout ),
	.dataf(!\F_ic_tag_rd_addr_nxt[3]~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_tag_rd_addr_nxt[4]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_tag_rd_addr_nxt[4]~13 .extended_lut = "off";
defparam \F_ic_tag_rd_addr_nxt[4]~13 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \F_ic_tag_rd_addr_nxt[4]~13 .shared_arith = "off";

dffeas \F_pc[7] (
	.clk(clk_clk),
	.d(\F_ic_tag_rd_addr_nxt[4]~13_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\F_pc[7]~q ),
	.prn(vcc));
defparam \F_pc[7] .is_wysiwyg = "true";
defparam \F_pc[7] .power_up = "low";

cyclonev_lcell_comb \Add3~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\F_pc[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~33_sumout ),
	.cout(\Add3~34 ),
	.shareout());
defparam \Add3~33 .extended_lut = "off";
defparam \Add3~33 .lut_mask = 64'h00000000000000FF;
defparam \Add3~33 .shared_arith = "off";

cyclonev_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[16] ),
	.datae(gnd),
	.dataf(!\Add3~33_sumout ),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout());
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~29 .shared_arith = "off";

dffeas \D_br_taken_waddr_partial[8] (
	.clk(clk_clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_br_taken_waddr_partial[8]~q ),
	.prn(vcc));
defparam \D_br_taken_waddr_partial[8] .is_wysiwyg = "true";
defparam \D_br_taken_waddr_partial[8] .power_up = "low";

cyclonev_lcell_comb \F_ic_tag_rd_addr_nxt[5]~14 (
	.dataa(!\D_pc[8]~q ),
	.datab(!\D_br_taken_waddr_partial[8]~q ),
	.datac(!\Add3~33_sumout ),
	.datad(!\D_iw[14]~q ),
	.datae(!\F_ic_tag_rd_addr_nxt[3]~0_combout ),
	.dataf(!\F_ic_tag_rd_addr_nxt[3]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_tag_rd_addr_nxt[5]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_tag_rd_addr_nxt[5]~14 .extended_lut = "off";
defparam \F_ic_tag_rd_addr_nxt[5]~14 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \F_ic_tag_rd_addr_nxt[5]~14 .shared_arith = "off";

dffeas \M_pc_plus_one[8] (
	.clk(clk_clk),
	.d(\Add7~25_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_pc_plus_one[8]~q ),
	.prn(vcc));
defparam \M_pc_plus_one[8] .is_wysiwyg = "true";
defparam \M_pc_plus_one[8] .power_up = "low";

dffeas \M_target_pcb[10] (
	.clk(clk_clk),
	.d(\E_src1[10]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_target_pcb[10]~q ),
	.prn(vcc));
defparam \M_target_pcb[10] .is_wysiwyg = "true";
defparam \M_target_pcb[10] .power_up = "low";

cyclonev_lcell_comb \A_pipe_flush_waddr_nxt~8 (
	.dataa(!\M_exc_any~combout ),
	.datab(!\M_pc_plus_one[8]~q ),
	.datac(!\M_ctrl_jmp_indirect~q ),
	.datad(!\M_target_pcb[10]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_pipe_flush_waddr_nxt~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_pipe_flush_waddr_nxt~8 .extended_lut = "off";
defparam \A_pipe_flush_waddr_nxt~8 .lut_mask = 64'hA3FFA3FFA3FFA3FF;
defparam \A_pipe_flush_waddr_nxt~8 .shared_arith = "off";

dffeas \A_pipe_flush_waddr[8] (
	.clk(clk_clk),
	.d(\A_pipe_flush_waddr_nxt~8_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\M_exc_break~0_combout ),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_pipe_flush_waddr[8]~q ),
	.prn(vcc));
defparam \A_pipe_flush_waddr[8] .is_wysiwyg = "true";
defparam \A_pipe_flush_waddr[8] .power_up = "low";

dffeas \D_pc_plus_one[8] (
	.clk(clk_clk),
	.d(\Add3~33_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_pc_plus_one[8]~q ),
	.prn(vcc));
defparam \D_pc_plus_one[8] .is_wysiwyg = "true";
defparam \D_pc_plus_one[8] .power_up = "low";

dffeas \E_extra_pc[8] (
	.clk(clk_clk),
	.d(\D_br_taken_waddr_partial[8]~q ),
	.asdata(\D_pc_plus_one[8]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_br_pred_not_taken~combout ),
	.ena(!\A_mem_stall~q ),
	.q(\E_extra_pc[8]~q ),
	.prn(vcc));
defparam \E_extra_pc[8] .is_wysiwyg = "true";
defparam \E_extra_pc[8] .power_up = "low";

dffeas \M_pipe_flush_waddr[8] (
	.clk(clk_clk),
	.d(\E_extra_pc[8]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_pipe_flush_waddr[8]~q ),
	.prn(vcc));
defparam \M_pipe_flush_waddr[8] .is_wysiwyg = "true";
defparam \M_pipe_flush_waddr[8] .power_up = "low";

cyclonev_lcell_comb \F_ic_tag_rd_addr_nxt[5]~15 (
	.dataa(!\F_ic_tag_rd_addr_nxt[5]~14_combout ),
	.datab(!\E_src1[10]~q ),
	.datac(!\A_pipe_flush_waddr[8]~q ),
	.datad(!\M_pipe_flush_waddr[8]~q ),
	.datae(!\F_ic_tag_rd_addr_nxt[3]~2_combout ),
	.dataf(!\F_ic_tag_rd_addr_nxt[3]~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_tag_rd_addr_nxt[5]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_tag_rd_addr_nxt[5]~15 .extended_lut = "off";
defparam \F_ic_tag_rd_addr_nxt[5]~15 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \F_ic_tag_rd_addr_nxt[5]~15 .shared_arith = "off";

dffeas \F_pc[8] (
	.clk(clk_clk),
	.d(\F_ic_tag_rd_addr_nxt[5]~15_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\F_pc[8]~q ),
	.prn(vcc));
defparam \F_pc[8] .is_wysiwyg = "true";
defparam \F_pc[8] .power_up = "low";

cyclonev_lcell_comb \Add3~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\F_pc[9]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~41_sumout ),
	.cout(\Add3~42 ),
	.shareout());
defparam \Add3~41 .extended_lut = "off";
defparam \Add3~41 .lut_mask = 64'h00000000000000FF;
defparam \Add3~41 .shared_arith = "off";

cyclonev_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[17] ),
	.datae(gnd),
	.dataf(!\Add3~41_sumout ),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~25 .shared_arith = "off";

dffeas \D_br_taken_waddr_partial[9] (
	.clk(clk_clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_br_taken_waddr_partial[9]~q ),
	.prn(vcc));
defparam \D_br_taken_waddr_partial[9] .is_wysiwyg = "true";
defparam \D_br_taken_waddr_partial[9] .power_up = "low";

cyclonev_lcell_comb \F_pc_nxt[9]~2 (
	.dataa(!\D_pc[9]~q ),
	.datab(!\D_br_taken_waddr_partial[9]~q ),
	.datac(!\Add3~41_sumout ),
	.datad(!\D_iw[15]~q ),
	.datae(!\F_ic_tag_rd_addr_nxt[3]~0_combout ),
	.dataf(!\F_ic_tag_rd_addr_nxt[3]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_pc_nxt[9]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_pc_nxt[9]~2 .extended_lut = "off";
defparam \F_pc_nxt[9]~2 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \F_pc_nxt[9]~2 .shared_arith = "off";

dffeas \M_target_pcb[11] (
	.clk(clk_clk),
	.d(\E_src1[11]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_target_pcb[11]~q ),
	.prn(vcc));
defparam \M_target_pcb[11] .is_wysiwyg = "true";
defparam \M_target_pcb[11] .power_up = "low";

cyclonev_lcell_comb \A_pipe_flush_waddr_nxt~10 (
	.dataa(!\M_exc_any~combout ),
	.datab(!\M_exc_break~0_combout ),
	.datac(!\M_pc_plus_one[9]~q ),
	.datad(!\M_ctrl_jmp_indirect~q ),
	.datae(!\M_target_pcb[11]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_pipe_flush_waddr_nxt~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_pipe_flush_waddr_nxt~10 .extended_lut = "off";
defparam \A_pipe_flush_waddr_nxt~10 .lut_mask = 64'hAF3FFFFFAF3FFFFF;
defparam \A_pipe_flush_waddr_nxt~10 .shared_arith = "off";

dffeas \A_pipe_flush_waddr[9] (
	.clk(clk_clk),
	.d(\A_pipe_flush_waddr_nxt~10_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_pipe_flush_waddr[9]~q ),
	.prn(vcc));
defparam \A_pipe_flush_waddr[9] .is_wysiwyg = "true";
defparam \A_pipe_flush_waddr[9] .power_up = "low";

dffeas \M_pipe_flush_waddr[9] (
	.clk(clk_clk),
	.d(\E_extra_pc[9]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_pipe_flush_waddr[9]~q ),
	.prn(vcc));
defparam \M_pipe_flush_waddr[9] .is_wysiwyg = "true";
defparam \M_pipe_flush_waddr[9] .power_up = "low";

cyclonev_lcell_comb \F_pc_nxt[9]~3 (
	.dataa(!\F_pc_nxt[9]~2_combout ),
	.datab(!\E_src1[11]~q ),
	.datac(!\A_pipe_flush_waddr[9]~q ),
	.datad(!\M_pipe_flush_waddr[9]~q ),
	.datae(!\F_ic_tag_rd_addr_nxt[3]~2_combout ),
	.dataf(!\F_ic_tag_rd_addr_nxt[3]~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_pc_nxt[9]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_pc_nxt[9]~3 .extended_lut = "off";
defparam \F_pc_nxt[9]~3 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \F_pc_nxt[9]~3 .shared_arith = "off";

dffeas \F_pc[9] (
	.clk(clk_clk),
	.d(\F_pc_nxt[9]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\F_pc[9]~q ),
	.prn(vcc));
defparam \F_pc[9] .is_wysiwyg = "true";
defparam \F_pc[9] .power_up = "low";

cyclonev_lcell_comb \Add3~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\F_pc[10]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~45_sumout ),
	.cout(\Add3~46 ),
	.shareout());
defparam \Add3~45 .extended_lut = "off";
defparam \Add3~45 .lut_mask = 64'h00000000000000FF;
defparam \Add3~45 .shared_arith = "off";

dffeas \D_pc_plus_one[10] (
	.clk(clk_clk),
	.d(\Add3~45_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_pc_plus_one[10]~q ),
	.prn(vcc));
defparam \D_pc_plus_one[10] .is_wysiwyg = "true";
defparam \D_pc_plus_one[10] .power_up = "low";

cyclonev_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(),
	.shareout());
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h0000000000000000;
defparam \Add0~41 .shared_arith = "off";

dffeas \D_br_taken_waddr_partial[10] (
	.clk(clk_clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_br_taken_waddr_partial[10]~q ),
	.prn(vcc));
defparam \D_br_taken_waddr_partial[10] .is_wysiwyg = "true";
defparam \D_br_taken_waddr_partial[10] .power_up = "low";

cyclonev_lcell_comb \Add1~22 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\D_br_taken_waddr_partial[10]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\Add1~22_cout ),
	.shareout());
defparam \Add1~22 .extended_lut = "off";
defparam \Add1~22 .lut_mask = 64'h00000000000000FF;
defparam \Add1~22 .shared_arith = "off";

cyclonev_lcell_comb \Add1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\D_pc_plus_one[10]~q ),
	.datae(gnd),
	.dataf(!\D_iw[18]~q ),
	.datag(gnd),
	.cin(\Add1~22_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~9_sumout ),
	.cout(\Add1~10 ),
	.shareout());
defparam \Add1~9 .extended_lut = "off";
defparam \Add1~9 .lut_mask = 64'h0000FF00000000FF;
defparam \Add1~9 .shared_arith = "off";

cyclonev_lcell_comb \F_pc_nxt[10]~4 (
	.dataa(!\D_pc[10]~q ),
	.datab(!\Add1~9_sumout ),
	.datac(!\Add3~45_sumout ),
	.datad(!\D_iw[16]~q ),
	.datae(!\F_ic_tag_rd_addr_nxt[3]~0_combout ),
	.dataf(!\F_ic_tag_rd_addr_nxt[3]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_pc_nxt[10]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_pc_nxt[10]~4 .extended_lut = "off";
defparam \F_pc_nxt[10]~4 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \F_pc_nxt[10]~4 .shared_arith = "off";

dffeas \M_target_pcb[12] (
	.clk(clk_clk),
	.d(\E_src1[12]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_target_pcb[12]~q ),
	.prn(vcc));
defparam \M_target_pcb[12] .is_wysiwyg = "true";
defparam \M_target_pcb[12] .power_up = "low";

cyclonev_lcell_comb \A_pipe_flush_waddr_nxt~11 (
	.dataa(!\M_exc_any~combout ),
	.datab(!\M_pc_plus_one[10]~q ),
	.datac(!\M_ctrl_jmp_indirect~q ),
	.datad(!\M_target_pcb[12]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_pipe_flush_waddr_nxt~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_pipe_flush_waddr_nxt~11 .extended_lut = "off";
defparam \A_pipe_flush_waddr_nxt~11 .lut_mask = 64'hA3FFA3FFA3FFA3FF;
defparam \A_pipe_flush_waddr_nxt~11 .shared_arith = "off";

dffeas \A_pipe_flush_waddr[10] (
	.clk(clk_clk),
	.d(\A_pipe_flush_waddr_nxt~11_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\M_exc_break~0_combout ),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_pipe_flush_waddr[10]~q ),
	.prn(vcc));
defparam \A_pipe_flush_waddr[10] .is_wysiwyg = "true";
defparam \A_pipe_flush_waddr[10] .power_up = "low";

dffeas \M_pipe_flush_waddr[10] (
	.clk(clk_clk),
	.d(\E_extra_pc[10]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_pipe_flush_waddr[10]~q ),
	.prn(vcc));
defparam \M_pipe_flush_waddr[10] .is_wysiwyg = "true";
defparam \M_pipe_flush_waddr[10] .power_up = "low";

cyclonev_lcell_comb \F_pc_nxt[10]~5 (
	.dataa(!\F_pc_nxt[10]~4_combout ),
	.datab(!\E_src1[12]~q ),
	.datac(!\A_pipe_flush_waddr[10]~q ),
	.datad(!\M_pipe_flush_waddr[10]~q ),
	.datae(!\F_ic_tag_rd_addr_nxt[3]~2_combout ),
	.dataf(!\F_ic_tag_rd_addr_nxt[3]~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_pc_nxt[10]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_pc_nxt[10]~5 .extended_lut = "off";
defparam \F_pc_nxt[10]~5 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \F_pc_nxt[10]~5 .shared_arith = "off";

dffeas \F_pc[10] (
	.clk(clk_clk),
	.d(\F_pc_nxt[10]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\F_pc[10]~q ),
	.prn(vcc));
defparam \F_pc[10] .is_wysiwyg = "true";
defparam \F_pc[10] .power_up = "low";

cyclonev_lcell_comb \Add3~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\F_pc[11]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~49_sumout ),
	.cout(\Add3~50 ),
	.shareout());
defparam \Add3~49 .extended_lut = "off";
defparam \Add3~49 .lut_mask = 64'h00000000000000FF;
defparam \Add3~49 .shared_arith = "off";

dffeas \D_pc_plus_one[11] (
	.clk(clk_clk),
	.d(\Add3~49_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_pc_plus_one[11]~q ),
	.prn(vcc));
defparam \D_pc_plus_one[11] .is_wysiwyg = "true";
defparam \D_pc_plus_one[11] .power_up = "low";

cyclonev_lcell_comb \Add1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\D_pc_plus_one[11]~q ),
	.datae(gnd),
	.dataf(!\D_iw[19]~q ),
	.datag(gnd),
	.cin(\Add1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~13_sumout ),
	.cout(\Add1~14 ),
	.shareout());
defparam \Add1~13 .extended_lut = "off";
defparam \Add1~13 .lut_mask = 64'h0000FF00000000FF;
defparam \Add1~13 .shared_arith = "off";

cyclonev_lcell_comb \F_pc_nxt[11]~6 (
	.dataa(!\D_pc[11]~q ),
	.datab(!\Add1~13_sumout ),
	.datac(!\Add3~49_sumout ),
	.datad(!\D_iw[17]~q ),
	.datae(!\F_ic_tag_rd_addr_nxt[3]~0_combout ),
	.dataf(!\F_ic_tag_rd_addr_nxt[3]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_pc_nxt[11]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_pc_nxt[11]~6 .extended_lut = "off";
defparam \F_pc_nxt[11]~6 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \F_pc_nxt[11]~6 .shared_arith = "off";

dffeas \M_target_pcb[13] (
	.clk(clk_clk),
	.d(\E_src1[13]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_target_pcb[13]~q ),
	.prn(vcc));
defparam \M_target_pcb[13] .is_wysiwyg = "true";
defparam \M_target_pcb[13] .power_up = "low";

cyclonev_lcell_comb \A_pipe_flush_waddr_nxt~12 (
	.dataa(!\M_exc_any~combout ),
	.datab(!\M_pc_plus_one[11]~q ),
	.datac(!\M_ctrl_jmp_indirect~q ),
	.datad(!\M_target_pcb[13]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_pipe_flush_waddr_nxt~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_pipe_flush_waddr_nxt~12 .extended_lut = "off";
defparam \A_pipe_flush_waddr_nxt~12 .lut_mask = 64'hA3FFA3FFA3FFA3FF;
defparam \A_pipe_flush_waddr_nxt~12 .shared_arith = "off";

dffeas \A_pipe_flush_waddr[11] (
	.clk(clk_clk),
	.d(\A_pipe_flush_waddr_nxt~12_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\M_exc_break~0_combout ),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_pipe_flush_waddr[11]~q ),
	.prn(vcc));
defparam \A_pipe_flush_waddr[11] .is_wysiwyg = "true";
defparam \A_pipe_flush_waddr[11] .power_up = "low";

dffeas \M_pipe_flush_waddr[11] (
	.clk(clk_clk),
	.d(\E_extra_pc[11]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_pipe_flush_waddr[11]~q ),
	.prn(vcc));
defparam \M_pipe_flush_waddr[11] .is_wysiwyg = "true";
defparam \M_pipe_flush_waddr[11] .power_up = "low";

cyclonev_lcell_comb \F_pc_nxt[11]~7 (
	.dataa(!\F_pc_nxt[11]~6_combout ),
	.datab(!\E_src1[13]~q ),
	.datac(!\A_pipe_flush_waddr[11]~q ),
	.datad(!\M_pipe_flush_waddr[11]~q ),
	.datae(!\F_ic_tag_rd_addr_nxt[3]~2_combout ),
	.dataf(!\F_ic_tag_rd_addr_nxt[3]~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_pc_nxt[11]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_pc_nxt[11]~7 .extended_lut = "off";
defparam \F_pc_nxt[11]~7 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \F_pc_nxt[11]~7 .shared_arith = "off";

dffeas \F_pc[11] (
	.clk(clk_clk),
	.d(\F_pc_nxt[11]~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\F_pc[11]~q ),
	.prn(vcc));
defparam \F_pc[11] .is_wysiwyg = "true";
defparam \F_pc[11] .power_up = "low";

cyclonev_lcell_comb \Add3~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\F_pc[12]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~53_sumout ),
	.cout(\Add3~54 ),
	.shareout());
defparam \Add3~53 .extended_lut = "off";
defparam \Add3~53 .lut_mask = 64'h00000000000000FF;
defparam \Add3~53 .shared_arith = "off";

dffeas \D_pc_plus_one[12] (
	.clk(clk_clk),
	.d(\Add3~53_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_pc_plus_one[12]~q ),
	.prn(vcc));
defparam \D_pc_plus_one[12] .is_wysiwyg = "true";
defparam \D_pc_plus_one[12] .power_up = "low";

cyclonev_lcell_comb \Add1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\D_pc_plus_one[12]~q ),
	.datae(gnd),
	.dataf(!\D_iw[20]~q ),
	.datag(gnd),
	.cin(\Add1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~17_sumout ),
	.cout(\Add1~18 ),
	.shareout());
defparam \Add1~17 .extended_lut = "off";
defparam \Add1~17 .lut_mask = 64'h0000FF00000000FF;
defparam \Add1~17 .shared_arith = "off";

cyclonev_lcell_comb \F_pc_nxt[12]~8 (
	.dataa(!\D_pc[12]~q ),
	.datab(!\Add1~17_sumout ),
	.datac(!\Add3~53_sumout ),
	.datad(!\D_iw[18]~q ),
	.datae(!\F_ic_tag_rd_addr_nxt[3]~0_combout ),
	.dataf(!\F_ic_tag_rd_addr_nxt[3]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_pc_nxt[12]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_pc_nxt[12]~8 .extended_lut = "off";
defparam \F_pc_nxt[12]~8 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \F_pc_nxt[12]~8 .shared_arith = "off";

dffeas \M_pc_plus_one[12] (
	.clk(clk_clk),
	.d(\Add7~53_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_pc_plus_one[12]~q ),
	.prn(vcc));
defparam \M_pc_plus_one[12] .is_wysiwyg = "true";
defparam \M_pc_plus_one[12] .power_up = "low";

dffeas \M_target_pcb[14] (
	.clk(clk_clk),
	.d(\E_src1[14]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_target_pcb[14]~q ),
	.prn(vcc));
defparam \M_target_pcb[14] .is_wysiwyg = "true";
defparam \M_target_pcb[14] .power_up = "low";

cyclonev_lcell_comb \A_pipe_flush_waddr_nxt~13 (
	.dataa(!\M_exc_any~combout ),
	.datab(!\M_pc_plus_one[12]~q ),
	.datac(!\M_ctrl_jmp_indirect~q ),
	.datad(!\M_target_pcb[14]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_pipe_flush_waddr_nxt~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_pipe_flush_waddr_nxt~13 .extended_lut = "off";
defparam \A_pipe_flush_waddr_nxt~13 .lut_mask = 64'hA3FFA3FFA3FFA3FF;
defparam \A_pipe_flush_waddr_nxt~13 .shared_arith = "off";

dffeas \A_pipe_flush_waddr[12] (
	.clk(clk_clk),
	.d(\A_pipe_flush_waddr_nxt~13_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\M_exc_break~0_combout ),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_pipe_flush_waddr[12]~q ),
	.prn(vcc));
defparam \A_pipe_flush_waddr[12] .is_wysiwyg = "true";
defparam \A_pipe_flush_waddr[12] .power_up = "low";

dffeas \E_extra_pc[12] (
	.clk(clk_clk),
	.d(\Add1~17_sumout ),
	.asdata(\D_pc_plus_one[12]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_br_pred_not_taken~combout ),
	.ena(!\A_mem_stall~q ),
	.q(\E_extra_pc[12]~q ),
	.prn(vcc));
defparam \E_extra_pc[12] .is_wysiwyg = "true";
defparam \E_extra_pc[12] .power_up = "low";

dffeas \M_pipe_flush_waddr[12] (
	.clk(clk_clk),
	.d(\E_extra_pc[12]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_pipe_flush_waddr[12]~q ),
	.prn(vcc));
defparam \M_pipe_flush_waddr[12] .is_wysiwyg = "true";
defparam \M_pipe_flush_waddr[12] .power_up = "low";

cyclonev_lcell_comb \F_pc_nxt[12]~9 (
	.dataa(!\F_pc_nxt[12]~8_combout ),
	.datab(!\E_src1[14]~q ),
	.datac(!\A_pipe_flush_waddr[12]~q ),
	.datad(!\M_pipe_flush_waddr[12]~q ),
	.datae(!\F_ic_tag_rd_addr_nxt[3]~2_combout ),
	.dataf(!\F_ic_tag_rd_addr_nxt[3]~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_pc_nxt[12]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_pc_nxt[12]~9 .extended_lut = "off";
defparam \F_pc_nxt[12]~9 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \F_pc_nxt[12]~9 .shared_arith = "off";

dffeas \F_pc[12] (
	.clk(clk_clk),
	.d(\F_pc_nxt[12]~9_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\F_pc[12]~q ),
	.prn(vcc));
defparam \F_pc[12] .is_wysiwyg = "true";
defparam \F_pc[12] .power_up = "low";

cyclonev_lcell_comb \Add3~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\F_pc[13]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~57_sumout ),
	.cout(\Add3~58 ),
	.shareout());
defparam \Add3~57 .extended_lut = "off";
defparam \Add3~57 .lut_mask = 64'h00000000000000FF;
defparam \Add3~57 .shared_arith = "off";

dffeas \D_pc_plus_one[13] (
	.clk(clk_clk),
	.d(\Add3~57_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_pc_plus_one[13]~q ),
	.prn(vcc));
defparam \D_pc_plus_one[13] .is_wysiwyg = "true";
defparam \D_pc_plus_one[13] .power_up = "low";

cyclonev_lcell_comb \Add1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\D_pc_plus_one[13]~q ),
	.datae(gnd),
	.dataf(!\D_iw[21]~q ),
	.datag(gnd),
	.cin(\Add1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~5_sumout ),
	.cout(\Add1~6 ),
	.shareout());
defparam \Add1~5 .extended_lut = "off";
defparam \Add1~5 .lut_mask = 64'h0000FF00000000FF;
defparam \Add1~5 .shared_arith = "off";

cyclonev_lcell_comb \F_pc_nxt[13]~10 (
	.dataa(!\D_pc[13]~q ),
	.datab(!\Add1~5_sumout ),
	.datac(!\Add3~57_sumout ),
	.datad(!\D_iw[19]~q ),
	.datae(!\F_ic_tag_rd_addr_nxt[3]~0_combout ),
	.dataf(!\F_ic_tag_rd_addr_nxt[3]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_pc_nxt[13]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_pc_nxt[13]~10 .extended_lut = "off";
defparam \F_pc_nxt[13]~10 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \F_pc_nxt[13]~10 .shared_arith = "off";

dffeas \M_target_pcb[15] (
	.clk(clk_clk),
	.d(\E_src1[15]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_target_pcb[15]~q ),
	.prn(vcc));
defparam \M_target_pcb[15] .is_wysiwyg = "true";
defparam \M_target_pcb[15] .power_up = "low";

cyclonev_lcell_comb \A_pipe_flush_waddr_nxt~14 (
	.dataa(!\M_exc_any~combout ),
	.datab(!\M_pc_plus_one[13]~q ),
	.datac(!\M_ctrl_jmp_indirect~q ),
	.datad(!\M_target_pcb[15]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_pipe_flush_waddr_nxt~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_pipe_flush_waddr_nxt~14 .extended_lut = "off";
defparam \A_pipe_flush_waddr_nxt~14 .lut_mask = 64'h53FF53FF53FF53FF;
defparam \A_pipe_flush_waddr_nxt~14 .shared_arith = "off";

dffeas \A_pipe_flush_waddr[13] (
	.clk(clk_clk),
	.d(\A_pipe_flush_waddr_nxt~14_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\M_exc_break~0_combout ),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_pipe_flush_waddr[13]~q ),
	.prn(vcc));
defparam \A_pipe_flush_waddr[13] .is_wysiwyg = "true";
defparam \A_pipe_flush_waddr[13] .power_up = "low";

cyclonev_lcell_comb \M_pipe_flush_waddr[13]~0 (
	.dataa(!\E_extra_pc[13]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_pipe_flush_waddr[13]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_pipe_flush_waddr[13]~0 .extended_lut = "off";
defparam \M_pipe_flush_waddr[13]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \M_pipe_flush_waddr[13]~0 .shared_arith = "off";

dffeas \M_pipe_flush_waddr[13] (
	.clk(clk_clk),
	.d(\M_pipe_flush_waddr[13]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_pipe_flush_waddr[13]~q ),
	.prn(vcc));
defparam \M_pipe_flush_waddr[13] .is_wysiwyg = "true";
defparam \M_pipe_flush_waddr[13] .power_up = "low";

cyclonev_lcell_comb \F_pc_nxt[13]~11 (
	.dataa(!\F_pc_nxt[13]~10_combout ),
	.datab(!\E_src1[15]~q ),
	.datac(!\A_pipe_flush_waddr[13]~q ),
	.datad(!\M_pipe_flush_waddr[13]~q ),
	.datae(!\F_ic_tag_rd_addr_nxt[3]~2_combout ),
	.dataf(!\F_ic_tag_rd_addr_nxt[3]~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_pc_nxt[13]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_pc_nxt[13]~11 .extended_lut = "off";
defparam \F_pc_nxt[13]~11 .lut_mask = 64'hFF7FFFFFFFFFFF7F;
defparam \F_pc_nxt[13]~11 .shared_arith = "off";

dffeas \F_pc[13] (
	.clk(clk_clk),
	.d(\F_pc_nxt[13]~11_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\F_pc[13]~q ),
	.prn(vcc));
defparam \F_pc[13] .is_wysiwyg = "true";
defparam \F_pc[13] .power_up = "low";

cyclonev_lcell_comb \Add3~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\F_pc[14]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~37_sumout ),
	.cout(),
	.shareout());
defparam \Add3~37 .extended_lut = "off";
defparam \Add3~37 .lut_mask = 64'h00000000000000FF;
defparam \Add3~37 .shared_arith = "off";

dffeas \D_pc_plus_one[14] (
	.clk(clk_clk),
	.d(\Add3~37_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_pc_plus_one[14]~q ),
	.prn(vcc));
defparam \D_pc_plus_one[14] .is_wysiwyg = "true";
defparam \D_pc_plus_one[14] .power_up = "low";

cyclonev_lcell_comb \Add1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\D_pc_plus_one[14]~q ),
	.datae(gnd),
	.dataf(!\D_iw[21]~q ),
	.datag(gnd),
	.cin(\Add1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~1_sumout ),
	.cout(),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h0000FF00000000FF;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \F_pc_nxt[14]~0 (
	.dataa(!\D_pc[14]~q ),
	.datab(!\Add1~1_sumout ),
	.datac(!\Add3~37_sumout ),
	.datad(!\D_iw[20]~q ),
	.datae(!\F_ic_tag_rd_addr_nxt[3]~0_combout ),
	.dataf(!\F_ic_tag_rd_addr_nxt[3]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_pc_nxt[14]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_pc_nxt[14]~0 .extended_lut = "off";
defparam \F_pc_nxt[14]~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \F_pc_nxt[14]~0 .shared_arith = "off";

dffeas \M_target_pcb[16] (
	.clk(clk_clk),
	.d(\E_src1[16]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_target_pcb[16]~q ),
	.prn(vcc));
defparam \M_target_pcb[16] .is_wysiwyg = "true";
defparam \M_target_pcb[16] .power_up = "low";

cyclonev_lcell_comb \A_pipe_flush_waddr_nxt~9 (
	.dataa(!\M_exc_any~combout ),
	.datab(!\M_exc_break~0_combout ),
	.datac(!\M_pc_plus_one[14]~q ),
	.datad(!\M_ctrl_jmp_indirect~q ),
	.datae(!\M_target_pcb[16]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_pipe_flush_waddr_nxt~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_pipe_flush_waddr_nxt~9 .extended_lut = "off";
defparam \A_pipe_flush_waddr_nxt~9 .lut_mask = 64'hAF3FFFFFAF3FFFFF;
defparam \A_pipe_flush_waddr_nxt~9 .shared_arith = "off";

dffeas \A_pipe_flush_waddr[14] (
	.clk(clk_clk),
	.d(\A_pipe_flush_waddr_nxt~9_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_pipe_flush_waddr[14]~q ),
	.prn(vcc));
defparam \A_pipe_flush_waddr[14] .is_wysiwyg = "true";
defparam \A_pipe_flush_waddr[14] .power_up = "low";

dffeas \M_pipe_flush_waddr[14] (
	.clk(clk_clk),
	.d(\E_extra_pc[14]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_pipe_flush_waddr[14]~q ),
	.prn(vcc));
defparam \M_pipe_flush_waddr[14] .is_wysiwyg = "true";
defparam \M_pipe_flush_waddr[14] .power_up = "low";

cyclonev_lcell_comb \F_pc_nxt[14]~1 (
	.dataa(!\F_pc_nxt[14]~0_combout ),
	.datab(!\E_src1[16]~q ),
	.datac(!\A_pipe_flush_waddr[14]~q ),
	.datad(!\M_pipe_flush_waddr[14]~q ),
	.datae(!\F_ic_tag_rd_addr_nxt[3]~2_combout ),
	.dataf(!\F_ic_tag_rd_addr_nxt[3]~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_pc_nxt[14]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_pc_nxt[14]~1 .extended_lut = "off";
defparam \F_pc_nxt[14]~1 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \F_pc_nxt[14]~1 .shared_arith = "off";

dffeas \F_pc[14] (
	.clk(clk_clk),
	.d(\F_pc_nxt[14]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\F_pc[14]~q ),
	.prn(vcc));
defparam \F_pc[14] .is_wysiwyg = "true";
defparam \F_pc[14] .power_up = "low";

cyclonev_lcell_comb \F_ic_hit~0 (
	.dataa(!\F_pc[9]~q ),
	.datab(!\first_nios2_system_cpu_cpu_ic_tag|the_altsyncram|auto_generated|q_b[0] ),
	.datac(!\F_pc[10]~q ),
	.datad(!\first_nios2_system_cpu_cpu_ic_tag|the_altsyncram|auto_generated|q_b[1] ),
	.datae(!\F_pc[11]~q ),
	.dataf(!\first_nios2_system_cpu_cpu_ic_tag|the_altsyncram|auto_generated|q_b[2] ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_hit~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_hit~0 .extended_lut = "off";
defparam \F_ic_hit~0 .lut_mask = 64'h6996966996696996;
defparam \F_ic_hit~0 .shared_arith = "off";

cyclonev_lcell_comb \F_ic_hit~1 (
	.dataa(!\F_pc[12]~q ),
	.datab(!\first_nios2_system_cpu_cpu_ic_tag|the_altsyncram|auto_generated|q_b[3] ),
	.datac(!\F_pc[13]~q ),
	.datad(!\first_nios2_system_cpu_cpu_ic_tag|the_altsyncram|auto_generated|q_b[4] ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_hit~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_hit~1 .extended_lut = "off";
defparam \F_ic_hit~1 .lut_mask = 64'h6996699669966996;
defparam \F_ic_hit~1 .shared_arith = "off";

cyclonev_lcell_comb F_ic_hit(
	.dataa(!\F_ic_valid~0_combout ),
	.datab(!\F_pc[14]~q ),
	.datac(!\first_nios2_system_cpu_cpu_ic_tag|the_altsyncram|auto_generated|q_b[5] ),
	.datad(!\F_ic_hit~0_combout ),
	.datae(!\F_ic_hit~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_hit~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam F_ic_hit.extended_lut = "off";
defparam F_ic_hit.lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam F_ic_hit.shared_arith = "off";

dffeas D_iw_valid(
	.clk(clk_clk),
	.d(\F_ic_hit~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_iw_valid~q ),
	.prn(vcc));
defparam D_iw_valid.is_wysiwyg = "true";
defparam D_iw_valid.power_up = "low";

cyclonev_lcell_comb \F_kill~0 (
	.dataa(!\M_pipe_flush~q ),
	.datab(!\E_valid_jmp_indirect~q ),
	.datac(!\D_iw_valid~q ),
	.datad(!\D_kill~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_kill~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_kill~0 .extended_lut = "off";
defparam \F_kill~0 .lut_mask = 64'hDFFFDFFFDFFFDFFF;
defparam \F_kill~0 .shared_arith = "off";

cyclonev_lcell_comb F_kill(
	.dataa(!\D_issue~q ),
	.datab(!\Equal95~4_combout ),
	.datac(!\Equal95~6_combout ),
	.datad(!\D_br_pred_taken~0_combout ),
	.datae(!\F_older_non_sequential~0_combout ),
	.dataf(!\F_kill~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_kill~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam F_kill.extended_lut = "off";
defparam F_kill.lut_mask = 64'hFFFFFFFF7FFFFFFF;
defparam F_kill.shared_arith = "off";

cyclonev_lcell_comb F_issue(
	.dataa(!\F_kill~combout ),
	.datab(!\F_ic_valid~0_combout ),
	.datac(!\F_pc[14]~q ),
	.datad(!\first_nios2_system_cpu_cpu_ic_tag|the_altsyncram|auto_generated|q_b[5] ),
	.datae(!\F_ic_hit~0_combout ),
	.dataf(!\F_ic_hit~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_issue~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam F_issue.extended_lut = "off";
defparam F_issue.lut_mask = 64'hBFFBFFFFFFFFFFFF;
defparam F_issue.shared_arith = "off";

dffeas D_issue(
	.clk(clk_clk),
	.d(\F_issue~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_issue~q ),
	.prn(vcc));
defparam D_issue.is_wysiwyg = "true";
defparam D_issue.power_up = "low";

cyclonev_lcell_comb \F_ic_tag_rd_addr_nxt[3]~0 (
	.dataa(!\D_issue~q ),
	.datab(!\D_ctrl_a_not_src~q ),
	.datac(!\D_iw_valid~q ),
	.datad(!\D_kill~q ),
	.datae(!\D_br_pred_taken~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_tag_rd_addr_nxt[3]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_tag_rd_addr_nxt[3]~0 .extended_lut = "off";
defparam \F_ic_tag_rd_addr_nxt[3]~0 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \F_ic_tag_rd_addr_nxt[3]~0 .shared_arith = "off";

cyclonev_lcell_comb \F_ic_tag_rd_addr_nxt[0]~4 (
	.dataa(!\D_pc[3]~q ),
	.datab(!\D_br_taken_waddr_partial[3]~q ),
	.datac(!\Add3~13_sumout ),
	.datad(!\D_iw[9]~q ),
	.datae(!\F_ic_tag_rd_addr_nxt[3]~0_combout ),
	.dataf(!\F_ic_tag_rd_addr_nxt[3]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_tag_rd_addr_nxt[0]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_tag_rd_addr_nxt[0]~4 .extended_lut = "off";
defparam \F_ic_tag_rd_addr_nxt[0]~4 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \F_ic_tag_rd_addr_nxt[0]~4 .shared_arith = "off";

dffeas \M_pc_plus_one[3] (
	.clk(clk_clk),
	.d(\Add7~9_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_pc_plus_one[3]~q ),
	.prn(vcc));
defparam \M_pc_plus_one[3] .is_wysiwyg = "true";
defparam \M_pc_plus_one[3] .power_up = "low";

dffeas \M_target_pcb[5] (
	.clk(clk_clk),
	.d(\E_src1[5]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_target_pcb[5]~q ),
	.prn(vcc));
defparam \M_target_pcb[5] .is_wysiwyg = "true";
defparam \M_target_pcb[5] .power_up = "low";

cyclonev_lcell_comb \A_pipe_flush_waddr_nxt~3 (
	.dataa(!\M_exc_any~combout ),
	.datab(!\M_pc_plus_one[3]~q ),
	.datac(!\M_ctrl_jmp_indirect~q ),
	.datad(!\M_target_pcb[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_pipe_flush_waddr_nxt~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_pipe_flush_waddr_nxt~3 .extended_lut = "off";
defparam \A_pipe_flush_waddr_nxt~3 .lut_mask = 64'h53FF53FF53FF53FF;
defparam \A_pipe_flush_waddr_nxt~3 .shared_arith = "off";

dffeas \A_pipe_flush_waddr[3] (
	.clk(clk_clk),
	.d(\A_pipe_flush_waddr_nxt~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_pipe_flush_waddr[3]~q ),
	.prn(vcc));
defparam \A_pipe_flush_waddr[3] .is_wysiwyg = "true";
defparam \A_pipe_flush_waddr[3] .power_up = "low";

dffeas \M_pipe_flush_waddr[3] (
	.clk(clk_clk),
	.d(\E_extra_pc[3]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_pipe_flush_waddr[3]~q ),
	.prn(vcc));
defparam \M_pipe_flush_waddr[3] .is_wysiwyg = "true";
defparam \M_pipe_flush_waddr[3] .power_up = "low";

cyclonev_lcell_comb \F_ic_tag_rd_addr_nxt[0]~5 (
	.dataa(!\F_ic_tag_rd_addr_nxt[0]~4_combout ),
	.datab(!\E_src1[5]~q ),
	.datac(!\A_pipe_flush_waddr[3]~q ),
	.datad(!\M_pipe_flush_waddr[3]~q ),
	.datae(!\F_ic_tag_rd_addr_nxt[3]~2_combout ),
	.dataf(!\F_ic_tag_rd_addr_nxt[3]~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_tag_rd_addr_nxt[0]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_tag_rd_addr_nxt[0]~5 .extended_lut = "off";
defparam \F_ic_tag_rd_addr_nxt[0]~5 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \F_ic_tag_rd_addr_nxt[0]~5 .shared_arith = "off";

dffeas \F_pc[3] (
	.clk(clk_clk),
	.d(\F_ic_tag_rd_addr_nxt[0]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\F_pc[3]~q ),
	.prn(vcc));
defparam \F_pc[3] .is_wysiwyg = "true";
defparam \F_pc[3] .power_up = "low";

dffeas \D_br_taken_waddr_partial[3] (
	.clk(clk_clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_br_taken_waddr_partial[3]~q ),
	.prn(vcc));
defparam \D_br_taken_waddr_partial[3] .is_wysiwyg = "true";
defparam \D_br_taken_waddr_partial[3] .power_up = "low";

dffeas \D_pc_plus_one[3] (
	.clk(clk_clk),
	.d(\Add3~13_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_pc_plus_one[3]~q ),
	.prn(vcc));
defparam \D_pc_plus_one[3] .is_wysiwyg = "true";
defparam \D_pc_plus_one[3] .power_up = "low";

dffeas \E_extra_pc[3] (
	.clk(clk_clk),
	.d(\D_br_taken_waddr_partial[3]~q ),
	.asdata(\D_pc_plus_one[3]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_br_pred_not_taken~combout ),
	.ena(!\A_mem_stall~q ),
	.q(\E_extra_pc[3]~q ),
	.prn(vcc));
defparam \E_extra_pc[3] .is_wysiwyg = "true";
defparam \E_extra_pc[3] .power_up = "low";

cyclonev_lcell_comb \E_alu_result[5] (
	.dataa(!\Add9~5_sumout ),
	.datab(!\E_ctrl_retaddr~q ),
	.datac(!\E_alu_result~0_combout ),
	.datad(!\E_alu_result~4_combout ),
	.datae(!\E_extra_pc[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[5]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[5] .extended_lut = "off";
defparam \E_alu_result[5] .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \E_alu_result[5] .shared_arith = "off";

dffeas \M_alu_result[5] (
	.clk(clk_clk),
	.d(\E_alu_result[5]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_alu_result[5]~q ),
	.prn(vcc));
defparam \M_alu_result[5] .is_wysiwyg = "true";
defparam \M_alu_result[5] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[5]~17 (
	.dataa(!\M_alu_result[5]~q ),
	.datab(!\A_wr_data_unfiltered[5]~7_combout ),
	.datac(!\first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[5] ),
	.datad(!\W_wr_data[5]~q ),
	.datae(!\E_src1[26]~0_combout ),
	.dataf(!\E_src1[26]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[5]~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[5]~17 .extended_lut = "off";
defparam \D_src1_reg[5]~17 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[5]~17 .shared_arith = "off";

dffeas \E_src1[5] (
	.clk(clk_clk),
	.d(\D_src1_reg[5]~17_combout ),
	.asdata(\E_alu_result[5]~combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\Equal303~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(!\A_mem_stall~q ),
	.q(\E_src1[5]~q ),
	.prn(vcc));
defparam \E_src1[5] .is_wysiwyg = "true";
defparam \E_src1[5] .power_up = "low";

cyclonev_lcell_comb \E_rot_step1[5]~14 (
	.dataa(!\E_src1[5]~q ),
	.datab(!\E_src1[4]~q ),
	.datac(!\E_src1[3]~q ),
	.datad(!\E_src1[2]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add10~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[5]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[5]~14 .extended_lut = "off";
defparam \E_rot_step1[5]~14 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[5]~14 .shared_arith = "off";

dffeas \M_rot_prestep2[5] (
	.clk(clk_clk),
	.d(\E_rot_step1[1]~9_combout ),
	.asdata(\E_rot_step1[5]~14_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add10~1_combout ),
	.ena(!\A_mem_stall~q ),
	.q(\M_rot_prestep2[5]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[5] .is_wysiwyg = "true";
defparam \M_rot_prestep2[5] .power_up = "low";

cyclonev_lcell_comb \M_rot[5]~5 (
	.dataa(!\M_rot_prestep2[5]~q ),
	.datab(!\M_rot_prestep2[29]~q ),
	.datac(!\M_rot_prestep2[21]~q ),
	.datad(!\M_rot_prestep2[13]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[5]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[5]~5 .extended_lut = "off";
defparam \M_rot[5]~5 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[5]~5 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~5 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_pass0~q ),
	.datac(!\M_rot_sel_fill0~q ),
	.datad(!\M_rot_mask[5]~q ),
	.datae(!\M_rot[5]~5_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~5 .extended_lut = "off";
defparam \A_shift_rot_result~5 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~5 .shared_arith = "off";

dffeas \A_shift_rot_result[5] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_shift_rot_result[5]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[5] .is_wysiwyg = "true";
defparam \A_shift_rot_result[5] .power_up = "low";

dffeas \A_inst_result[5] (
	.clk(clk_clk),
	.d(\M_pc_plus_one[3]~q ),
	.asdata(\M_alu_result[5]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\A_inst_result[9]~0_combout ),
	.sload(!\M_exc_any~combout ),
	.ena(!\A_mem_stall~q ),
	.q(\A_inst_result[5]~q ),
	.prn(vcc));
defparam \A_inst_result[5] .is_wysiwyg = "true";
defparam \A_inst_result[5] .power_up = "low";

dffeas \A_mul_cell_p1[5] (
	.clk(clk_clk),
	.d(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[5]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_mul_cell_p1[5]~q ),
	.prn(vcc));
defparam \A_mul_cell_p1[5] .is_wysiwyg = "true";
defparam \A_mul_cell_p1[5] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[5]~7 (
	.dataa(!\A_slow_inst_result[5]~q ),
	.datab(!\A_shift_rot_result[5]~q ),
	.datac(!\A_inst_result[5]~q ),
	.datad(!\A_mul_cell_p1[5]~q ),
	.datae(!\A_wr_data_unfiltered[15]~0_combout ),
	.dataf(!\A_wr_data_unfiltered[15]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[5]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[5]~7 .extended_lut = "off";
defparam \A_wr_data_unfiltered[5]~7 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_wr_data_unfiltered[5]~7 .shared_arith = "off";

dffeas \W_wr_data[5] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[5]~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[5]~q ),
	.prn(vcc));
defparam \W_wr_data[5] .is_wysiwyg = "true";
defparam \W_wr_data[5] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[5]~20 (
	.dataa(!\D_src2_reg[0]~7_combout ),
	.datab(!\D_src2_reg[0]~8_combout ),
	.datac(!\W_wr_data[5]~q ),
	.datad(!\A_wr_data_unfiltered[5]~7_combout ),
	.datae(!\M_alu_result[5]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[5]~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[5]~20 .extended_lut = "off";
defparam \D_src2_reg[5]~20 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \D_src2_reg[5]~20 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[5]~21 (
	.dataa(!\D_src2_reg[0]~4_combout ),
	.datab(!\D_src2_reg[0]~5_combout ),
	.datac(!\D_src2_reg[5]~20_combout ),
	.datad(!\E_alu_result[5]~combout ),
	.datae(!\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[5] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[5]~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[5]~21 .extended_lut = "off";
defparam \D_src2_reg[5]~21 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \D_src2_reg[5]~21 .shared_arith = "off";

dffeas \E_src2[5] (
	.clk(clk_clk),
	.d(\D_iw[11]~q ),
	.asdata(\D_src2_reg[5]~21_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src2[5]~2_combout ),
	.sload(!\D_ctrl_src2_choose_imm~q ),
	.ena(!\A_mem_stall~q ),
	.q(\E_src2[5]~q ),
	.prn(vcc));
defparam \E_src2[5] .is_wysiwyg = "true";
defparam \E_src2[5] .power_up = "low";

cyclonev_lcell_comb \Add9~49 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[6]~q ),
	.datae(gnd),
	.dataf(!\E_src1[6]~q ),
	.datag(gnd),
	.cin(\Add9~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~49_sumout ),
	.cout(\Add9~50 ),
	.shareout());
defparam \Add9~49 .extended_lut = "off";
defparam \Add9~49 .lut_mask = 64'h0000FF00000055AA;
defparam \Add9~49 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result~6 (
	.dataa(!\E_src2[7]~q ),
	.datab(!\E_src1[7]~q ),
	.datac(!\E_logic_op[1]~q ),
	.datad(!\E_logic_op[0]~q ),
	.datae(!\E_ctrl_logic~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result~6 .extended_lut = "off";
defparam \E_alu_result~6 .lut_mask = 64'h6996FFFF6996FFFF;
defparam \E_alu_result~6 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[7] (
	.dataa(!\Add9~45_sumout ),
	.datab(!\E_ctrl_retaddr~q ),
	.datac(!\E_alu_result~0_combout ),
	.datad(!\E_alu_result~6_combout ),
	.datae(!\E_extra_pc[5]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[7]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[7] .extended_lut = "off";
defparam \E_alu_result[7] .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \E_alu_result[7] .shared_arith = "off";

dffeas \M_alu_result[7] (
	.clk(clk_clk),
	.d(\E_alu_result[7]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_alu_result[7]~q ),
	.prn(vcc));
defparam \M_alu_result[7] .is_wysiwyg = "true";
defparam \M_alu_result[7] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[7]~8 (
	.dataa(!\M_alu_result[7]~q ),
	.datab(!\A_wr_data_unfiltered[7]~9_combout ),
	.datac(!\first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[7] ),
	.datad(!\W_wr_data[7]~q ),
	.datae(!\E_src1[26]~0_combout ),
	.dataf(!\E_src1[26]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[7]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[7]~8 .extended_lut = "off";
defparam \D_src1_reg[7]~8 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[7]~8 .shared_arith = "off";

dffeas \E_src1[7] (
	.clk(clk_clk),
	.d(\D_src1_reg[7]~8_combout ),
	.asdata(\E_alu_result[7]~combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\Equal303~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(!\A_mem_stall~q ),
	.q(\E_src1[7]~q ),
	.prn(vcc));
defparam \E_src1[7] .is_wysiwyg = "true";
defparam \E_src1[7] .power_up = "low";

cyclonev_lcell_comb \E_rot_step1[7]~30 (
	.dataa(!\E_src1[7]~q ),
	.datab(!\E_src1[6]~q ),
	.datac(!\E_src1[5]~q ),
	.datad(!\E_src1[4]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add10~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[7]~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[7]~30 .extended_lut = "off";
defparam \E_rot_step1[7]~30 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[7]~30 .shared_arith = "off";

dffeas \M_rot_prestep2[7] (
	.clk(clk_clk),
	.d(\E_rot_step1[3]~25_combout ),
	.asdata(\E_rot_step1[7]~30_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add10~1_combout ),
	.ena(!\A_mem_stall~q ),
	.q(\M_rot_prestep2[7]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[7] .is_wysiwyg = "true";
defparam \M_rot_prestep2[7] .power_up = "low";

cyclonev_lcell_comb \M_rot[7]~7 (
	.dataa(!\M_rot_prestep2[7]~q ),
	.datab(!\M_rot_prestep2[31]~q ),
	.datac(!\M_rot_prestep2[23]~q ),
	.datad(!\M_rot_prestep2[15]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[7]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[7]~7 .extended_lut = "off";
defparam \M_rot[7]~7 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[7]~7 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~7 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_pass0~q ),
	.datac(!\M_rot_sel_fill0~q ),
	.datad(!\M_rot_mask[7]~q ),
	.datae(!\M_rot[7]~7_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~7 .extended_lut = "off";
defparam \A_shift_rot_result~7 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~7 .shared_arith = "off";

dffeas \A_shift_rot_result[7] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_shift_rot_result[7]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[7] .is_wysiwyg = "true";
defparam \A_shift_rot_result[7] .power_up = "low";

dffeas \A_inst_result[7] (
	.clk(clk_clk),
	.d(\M_pc_plus_one[5]~q ),
	.asdata(\M_alu_result[7]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\A_inst_result[9]~0_combout ),
	.sload(!\M_exc_any~combout ),
	.ena(!\A_mem_stall~q ),
	.q(\A_inst_result[7]~q ),
	.prn(vcc));
defparam \A_inst_result[7] .is_wysiwyg = "true";
defparam \A_inst_result[7] .power_up = "low";

dffeas \A_mul_cell_p1[7] (
	.clk(clk_clk),
	.d(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[7]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_mul_cell_p1[7]~q ),
	.prn(vcc));
defparam \A_mul_cell_p1[7] .is_wysiwyg = "true";
defparam \A_mul_cell_p1[7] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[7]~9 (
	.dataa(!\A_slow_inst_result[7]~q ),
	.datab(!\A_shift_rot_result[7]~q ),
	.datac(!\A_inst_result[7]~q ),
	.datad(!\A_mul_cell_p1[7]~q ),
	.datae(!\A_wr_data_unfiltered[15]~0_combout ),
	.dataf(!\A_wr_data_unfiltered[15]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[7]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[7]~9 .extended_lut = "off";
defparam \A_wr_data_unfiltered[7]~9 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_wr_data_unfiltered[7]~9 .shared_arith = "off";

dffeas \W_wr_data[7] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[7]~9_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[7]~q ),
	.prn(vcc));
defparam \W_wr_data[7] .is_wysiwyg = "true";
defparam \W_wr_data[7] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[7]~24 (
	.dataa(!\D_src2_reg[0]~7_combout ),
	.datab(!\D_src2_reg[0]~8_combout ),
	.datac(!\W_wr_data[7]~q ),
	.datad(!\A_wr_data_unfiltered[7]~9_combout ),
	.datae(!\M_alu_result[7]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[7]~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[7]~24 .extended_lut = "off";
defparam \D_src2_reg[7]~24 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \D_src2_reg[7]~24 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[7]~25 (
	.dataa(!\D_src2_reg[0]~4_combout ),
	.datab(!\D_src2_reg[0]~5_combout ),
	.datac(!\D_src2_reg[7]~24_combout ),
	.datad(!\E_alu_result[7]~combout ),
	.datae(!\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[7] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[7]~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[7]~25 .extended_lut = "off";
defparam \D_src2_reg[7]~25 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \D_src2_reg[7]~25 .shared_arith = "off";

dffeas \E_src2[7] (
	.clk(clk_clk),
	.d(\D_iw[13]~q ),
	.asdata(\D_src2_reg[7]~25_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src2[5]~2_combout ),
	.sload(!\D_ctrl_src2_choose_imm~q ),
	.ena(!\A_mem_stall~q ),
	.q(\E_src2[7]~q ),
	.prn(vcc));
defparam \E_src2[7] .is_wysiwyg = "true";
defparam \E_src2[7] .power_up = "low";

cyclonev_lcell_comb \Equal316~3 (
	.dataa(!\E_src2[7]~q ),
	.datab(!\E_src1[7]~q ),
	.datac(!\E_src2[21]~q ),
	.datad(!\E_src1[21]~q ),
	.datae(!\E_logic_op[1]~q ),
	.dataf(!\E_logic_op[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal316~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal316~3 .extended_lut = "off";
defparam \Equal316~3 .lut_mask = 64'h6996966996696996;
defparam \Equal316~3 .shared_arith = "off";

cyclonev_lcell_comb \Equal316~4 (
	.dataa(!\E_src2[11]~q ),
	.datab(!\E_src1[11]~q ),
	.datac(!\E_src2[28]~q ),
	.datad(!\E_src1[28]~q ),
	.datae(!\E_logic_op[1]~q ),
	.dataf(!\E_logic_op[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal316~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal316~4 .extended_lut = "off";
defparam \Equal316~4 .lut_mask = 64'h6996966996696996;
defparam \Equal316~4 .shared_arith = "off";

cyclonev_lcell_comb \Equal316~5 (
	.dataa(!\E_src2[10]~q ),
	.datab(!\E_src1[10]~q ),
	.datac(!\E_src2[27]~q ),
	.datad(!\E_src1[27]~q ),
	.datae(!\E_logic_op[1]~q ),
	.dataf(!\E_logic_op[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal316~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal316~5 .extended_lut = "off";
defparam \Equal316~5 .lut_mask = 64'h6996966996696996;
defparam \Equal316~5 .shared_arith = "off";

cyclonev_lcell_comb \Equal316~6 (
	.dataa(!\E_src2[8]~q ),
	.datab(!\E_src1[8]~q ),
	.datac(!\E_src2[9]~q ),
	.datad(!\E_src1[9]~q ),
	.datae(!\E_logic_op[1]~q ),
	.dataf(!\E_logic_op[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal316~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal316~6 .extended_lut = "off";
defparam \Equal316~6 .lut_mask = 64'h6996966996696996;
defparam \Equal316~6 .shared_arith = "off";

cyclonev_lcell_comb \Equal316~7 (
	.dataa(!\E_src2[4]~q ),
	.datab(!\E_src1[4]~q ),
	.datac(!\E_src2[5]~q ),
	.datad(!\E_src1[5]~q ),
	.datae(!\E_logic_op[1]~q ),
	.dataf(!\E_logic_op[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal316~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal316~7 .extended_lut = "off";
defparam \Equal316~7 .lut_mask = 64'h6996966996696996;
defparam \Equal316~7 .shared_arith = "off";

cyclonev_lcell_comb \Equal316~8 (
	.dataa(!\E_src2[6]~q ),
	.datab(!\E_src1[6]~q ),
	.datac(!\E_src2[26]~q ),
	.datad(!\E_src1[26]~q ),
	.datae(!\E_logic_op[1]~q ),
	.dataf(!\E_logic_op[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal316~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal316~8 .extended_lut = "off";
defparam \Equal316~8 .lut_mask = 64'h6996966996696996;
defparam \Equal316~8 .shared_arith = "off";

cyclonev_lcell_comb \Equal316~9 (
	.dataa(!\Equal316~3_combout ),
	.datab(!\Equal316~4_combout ),
	.datac(!\Equal316~5_combout ),
	.datad(!\Equal316~6_combout ),
	.datae(!\Equal316~7_combout ),
	.dataf(!\Equal316~8_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal316~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal316~9 .extended_lut = "off";
defparam \Equal316~9 .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \Equal316~9 .shared_arith = "off";

cyclonev_lcell_comb \Equal316~10 (
	.dataa(!\E_src2[20]~q ),
	.datab(!\E_src1[20]~q ),
	.datac(!\E_src2[19]~q ),
	.datad(!\E_src1[19]~q ),
	.datae(!\E_logic_op[1]~q ),
	.dataf(!\E_logic_op[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal316~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal316~10 .extended_lut = "off";
defparam \Equal316~10 .lut_mask = 64'h6996966996696996;
defparam \Equal316~10 .shared_arith = "off";

cyclonev_lcell_comb \Equal316~11 (
	.dataa(!\E_src2[1]~q ),
	.datab(!\E_src1[1]~q ),
	.datac(!\E_src2[18]~q ),
	.datad(!\E_src1[18]~q ),
	.datae(!\E_logic_op[1]~q ),
	.dataf(!\E_logic_op[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal316~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal316~11 .extended_lut = "off";
defparam \Equal316~11 .lut_mask = 64'h6996966996696996;
defparam \Equal316~11 .shared_arith = "off";

cyclonev_lcell_comb \Equal316~12 (
	.dataa(!\E_src2[16]~q ),
	.datab(!\E_src1[16]~q ),
	.datac(!\E_src2[15]~q ),
	.datad(!\E_src1[15]~q ),
	.datae(!\E_logic_op[1]~q ),
	.dataf(!\E_logic_op[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal316~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal316~12 .extended_lut = "off";
defparam \Equal316~12 .lut_mask = 64'h6996966996696996;
defparam \Equal316~12 .shared_arith = "off";

cyclonev_lcell_comb \Equal316~13 (
	.dataa(!\E_src2[12]~q ),
	.datab(!\E_src1[12]~q ),
	.datac(!\E_src2[13]~q ),
	.datad(!\E_src1[13]~q ),
	.datae(!\E_logic_op[1]~q ),
	.dataf(!\E_logic_op[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal316~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal316~13 .extended_lut = "off";
defparam \Equal316~13 .lut_mask = 64'h6996966996696996;
defparam \Equal316~13 .shared_arith = "off";

cyclonev_lcell_comb \Equal316~14 (
	.dataa(!\E_src2[14]~q ),
	.datab(!\E_src1[14]~q ),
	.datac(!\E_src2[29]~q ),
	.datad(!\E_src1[29]~q ),
	.datae(!\E_logic_op[1]~q ),
	.dataf(!\E_logic_op[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal316~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal316~14 .extended_lut = "off";
defparam \Equal316~14 .lut_mask = 64'h6996966996696996;
defparam \Equal316~14 .shared_arith = "off";

cyclonev_lcell_comb \Equal316~15 (
	.dataa(!\E_logic_result[17]~4_combout ),
	.datab(!\E_logic_result[30]~5_combout ),
	.datac(!\Equal316~11_combout ),
	.datad(!\Equal316~12_combout ),
	.datae(!\Equal316~13_combout ),
	.dataf(!\Equal316~14_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal316~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal316~15 .extended_lut = "off";
defparam \Equal316~15 .lut_mask = 64'hEFFFFFFFFFFFFFFF;
defparam \Equal316~15 .shared_arith = "off";

dffeas \E_compare_op[1] (
	.clk(clk_clk),
	.d(\D_logic_op_raw[1]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_compare_op[1]~q ),
	.prn(vcc));
defparam \E_compare_op[1] .is_wysiwyg = "true";
defparam \E_compare_op[1] .power_up = "low";

cyclonev_lcell_comb \E_br_result~0 (
	.dataa(!\E_compare_op[0]~q ),
	.datab(!\Equal316~2_combout ),
	.datac(!\Equal316~9_combout ),
	.datad(!\Equal316~10_combout ),
	.datae(!\Equal316~15_combout ),
	.dataf(!\E_compare_op[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_br_result~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_br_result~0 .extended_lut = "off";
defparam \E_br_result~0 .lut_mask = 64'hFFFFFFFF7DD7D77D;
defparam \E_br_result~0 .shared_arith = "off";

cyclonev_lcell_comb \E_br_result~1 (
	.dataa(!\E_compare_op[0]~q ),
	.datab(!\Equal316~2_combout ),
	.datac(!\Equal316~9_combout ),
	.datad(!\Equal316~10_combout ),
	.datae(!\Equal316~15_combout ),
	.dataf(!\E_compare_op[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_br_result~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_br_result~1 .extended_lut = "off";
defparam \E_br_result~1 .lut_mask = 64'hBEEBEBBEFFFFFFFF;
defparam \E_br_result~1 .shared_arith = "off";

cyclonev_lcell_comb \E_logic_result[0]~6 (
	.dataa(!\E_src2[0]~q ),
	.datab(!\E_src1[0]~q ),
	.datac(!\E_logic_op[1]~q ),
	.datad(!\E_logic_op[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[0]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[0]~6 .extended_lut = "off";
defparam \E_logic_result[0]~6 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[0]~6 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[0]~1 (
	.dataa(!\E_logic_result[0]~6_combout ),
	.datab(!\E_ctrl_logic~q ),
	.datac(!\Add9~65_sumout ),
	.datad(!\E_alu_result~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[0]~1 .extended_lut = "off";
defparam \E_alu_result[0]~1 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \E_alu_result[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[0] (
	.dataa(!\E_ctrl_cmp~q ),
	.datab(!\Add9~61_sumout ),
	.datac(!\E_br_result~0_combout ),
	.datad(!\E_br_result~1_combout ),
	.datae(!\E_alu_result[0]~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[0]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[0] .extended_lut = "off";
defparam \E_alu_result[0] .lut_mask = 64'h47FFFFFF47FFFFFF;
defparam \E_alu_result[0] .shared_arith = "off";

dffeas \M_alu_result[0] (
	.clk(clk_clk),
	.d(\E_alu_result[0]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_alu_result[0]~q ),
	.prn(vcc));
defparam \M_alu_result[0] .is_wysiwyg = "true";
defparam \M_alu_result[0] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[0]~4 (
	.dataa(!\M_alu_result[0]~q ),
	.datab(!\A_wr_data_unfiltered[0]~2_combout ),
	.datac(!\first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[0] ),
	.datad(!\W_wr_data[0]~q ),
	.datae(!\E_src1[26]~0_combout ),
	.dataf(!\E_src1[26]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[0]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[0]~4 .extended_lut = "off";
defparam \D_src1_reg[0]~4 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[0]~4 .shared_arith = "off";

dffeas \E_src1[0] (
	.clk(clk_clk),
	.d(\D_src1_reg[0]~4_combout ),
	.asdata(\E_alu_result[0]~combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\Equal303~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(!\A_mem_stall~q ),
	.q(\E_src1[0]~q ),
	.prn(vcc));
defparam \E_src1[0] .is_wysiwyg = "true";
defparam \E_src1[0] .power_up = "low";

cyclonev_lcell_comb \E_rot_step1[2]~17 (
	.dataa(!\E_src1[2]~q ),
	.datab(!\E_src1[1]~q ),
	.datac(!\E_src1[0]~q ),
	.datad(!\E_src1[31]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add10~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[2]~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[2]~17 .extended_lut = "off";
defparam \E_rot_step1[2]~17 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[2]~17 .shared_arith = "off";

dffeas \M_rot_prestep2[6] (
	.clk(clk_clk),
	.d(\E_rot_step1[2]~17_combout ),
	.asdata(\E_rot_step1[6]~22_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add10~1_combout ),
	.ena(!\A_mem_stall~q ),
	.q(\M_rot_prestep2[6]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[6] .is_wysiwyg = "true";
defparam \M_rot_prestep2[6] .power_up = "low";

cyclonev_lcell_comb \E_rot_step1[26]~19 (
	.dataa(!\E_src1[26]~q ),
	.datab(!\E_src1[25]~q ),
	.datac(!\E_src1[24]~q ),
	.datad(!\E_src1[23]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add10~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[26]~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[26]~19 .extended_lut = "off";
defparam \E_rot_step1[26]~19 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[26]~19 .shared_arith = "off";

dffeas \M_rot_prestep2[30] (
	.clk(clk_clk),
	.d(\E_rot_step1[26]~19_combout ),
	.asdata(\E_rot_step1[30]~16_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add10~1_combout ),
	.ena(!\A_mem_stall~q ),
	.q(\M_rot_prestep2[30]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[30] .is_wysiwyg = "true";
defparam \M_rot_prestep2[30] .power_up = "low";

cyclonev_lcell_comb \M_rot[6]~6 (
	.dataa(!\M_rot_prestep2[6]~q ),
	.datab(!\M_rot_prestep2[30]~q ),
	.datac(!\M_rot_prestep2[22]~q ),
	.datad(!\M_rot_prestep2[14]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[6]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[6]~6 .extended_lut = "off";
defparam \M_rot[6]~6 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[6]~6 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~6 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_pass0~q ),
	.datac(!\M_rot_sel_fill0~q ),
	.datad(!\M_rot_mask[6]~q ),
	.datae(!\M_rot[6]~6_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~6 .extended_lut = "off";
defparam \A_shift_rot_result~6 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~6 .shared_arith = "off";

dffeas \A_shift_rot_result[6] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_shift_rot_result[6]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[6] .is_wysiwyg = "true";
defparam \A_shift_rot_result[6] .power_up = "low";

dffeas \A_inst_result[6] (
	.clk(clk_clk),
	.d(\M_pc_plus_one[4]~q ),
	.asdata(\M_alu_result[6]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\A_inst_result[9]~0_combout ),
	.sload(!\M_exc_any~combout ),
	.ena(!\A_mem_stall~q ),
	.q(\A_inst_result[6]~q ),
	.prn(vcc));
defparam \A_inst_result[6] .is_wysiwyg = "true";
defparam \A_inst_result[6] .power_up = "low";

dffeas \A_mul_cell_p1[6] (
	.clk(clk_clk),
	.d(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[6]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_mul_cell_p1[6]~q ),
	.prn(vcc));
defparam \A_mul_cell_p1[6] .is_wysiwyg = "true";
defparam \A_mul_cell_p1[6] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[6]~8 (
	.dataa(!\A_slow_inst_result[6]~q ),
	.datab(!\A_shift_rot_result[6]~q ),
	.datac(!\A_inst_result[6]~q ),
	.datad(!\A_mul_cell_p1[6]~q ),
	.datae(!\A_wr_data_unfiltered[15]~0_combout ),
	.dataf(!\A_wr_data_unfiltered[15]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[6]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[6]~8 .extended_lut = "off";
defparam \A_wr_data_unfiltered[6]~8 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_wr_data_unfiltered[6]~8 .shared_arith = "off";

dffeas \W_wr_data[6] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[6]~8_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[6]~q ),
	.prn(vcc));
defparam \W_wr_data[6] .is_wysiwyg = "true";
defparam \W_wr_data[6] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[6]~22 (
	.dataa(!\D_src2_reg[0]~7_combout ),
	.datab(!\D_src2_reg[0]~8_combout ),
	.datac(!\W_wr_data[6]~q ),
	.datad(!\A_wr_data_unfiltered[6]~8_combout ),
	.datae(!\M_alu_result[6]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[6]~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[6]~22 .extended_lut = "off";
defparam \D_src2_reg[6]~22 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \D_src2_reg[6]~22 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[6]~23 (
	.dataa(!\D_src2_reg[0]~4_combout ),
	.datab(!\D_src2_reg[0]~5_combout ),
	.datac(!\D_src2_reg[6]~22_combout ),
	.datad(!\E_alu_result[6]~combout ),
	.datae(!\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[6] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[6]~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[6]~23 .extended_lut = "off";
defparam \D_src2_reg[6]~23 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \D_src2_reg[6]~23 .shared_arith = "off";

dffeas \E_src2[6] (
	.clk(clk_clk),
	.d(\D_iw[12]~q ),
	.asdata(\D_src2_reg[6]~23_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src2[5]~2_combout ),
	.sload(!\D_ctrl_src2_choose_imm~q ),
	.ena(!\A_mem_stall~q ),
	.q(\E_src2[6]~q ),
	.prn(vcc));
defparam \E_src2[6] .is_wysiwyg = "true";
defparam \E_src2[6] .power_up = "low";

cyclonev_lcell_comb \E_alu_result~5 (
	.dataa(!\E_src2[6]~q ),
	.datab(!\E_src1[6]~q ),
	.datac(!\E_logic_op[1]~q ),
	.datad(!\E_logic_op[0]~q ),
	.datae(!\E_ctrl_logic~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result~5 .extended_lut = "off";
defparam \E_alu_result~5 .lut_mask = 64'h6996FFFF6996FFFF;
defparam \E_alu_result~5 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[6] (
	.dataa(!\Add9~49_sumout ),
	.datab(!\E_ctrl_retaddr~q ),
	.datac(!\E_alu_result~0_combout ),
	.datad(!\E_alu_result~5_combout ),
	.datae(!\E_extra_pc[4]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[6]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[6] .extended_lut = "off";
defparam \E_alu_result[6] .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \E_alu_result[6] .shared_arith = "off";

dffeas \M_alu_result[6] (
	.clk(clk_clk),
	.d(\E_alu_result[6]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_alu_result[6]~q ),
	.prn(vcc));
defparam \M_alu_result[6] .is_wysiwyg = "true";
defparam \M_alu_result[6] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[6]~18 (
	.dataa(!\M_alu_result[6]~q ),
	.datab(!\A_wr_data_unfiltered[6]~8_combout ),
	.datac(!\first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[6] ),
	.datad(!\W_wr_data[6]~q ),
	.datae(!\E_src1[26]~0_combout ),
	.dataf(!\E_src1[26]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[6]~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[6]~18 .extended_lut = "off";
defparam \D_src1_reg[6]~18 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[6]~18 .shared_arith = "off";

dffeas \E_src1[6] (
	.clk(clk_clk),
	.d(\D_src1_reg[6]~18_combout ),
	.asdata(\E_alu_result[6]~combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\Equal303~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(!\A_mem_stall~q ),
	.q(\E_src1[6]~q ),
	.prn(vcc));
defparam \E_src1[6] .is_wysiwyg = "true";
defparam \E_src1[6] .power_up = "low";

cyclonev_lcell_comb \E_rot_step1[6]~22 (
	.dataa(!\E_src1[6]~q ),
	.datab(!\E_src1[5]~q ),
	.datac(!\E_src1[4]~q ),
	.datad(!\E_src1[3]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add10~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[6]~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[6]~22 .extended_lut = "off";
defparam \E_rot_step1[6]~22 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[6]~22 .shared_arith = "off";

dffeas \M_rot_prestep2[10] (
	.clk(clk_clk),
	.d(\E_rot_step1[6]~22_combout ),
	.asdata(\E_rot_step1[10]~23_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add10~1_combout ),
	.ena(!\A_mem_stall~q ),
	.q(\M_rot_prestep2[10]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[10] .is_wysiwyg = "true";
defparam \M_rot_prestep2[10] .power_up = "low";

cyclonev_lcell_comb \E_rot_step1[22]~18 (
	.dataa(!\E_src1[22]~q ),
	.datab(!\E_src1[21]~q ),
	.datac(!\E_src1[20]~q ),
	.datad(!\E_src1[19]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add10~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[22]~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[22]~18 .extended_lut = "off";
defparam \E_rot_step1[22]~18 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[22]~18 .shared_arith = "off";

dffeas \M_rot_prestep2[26] (
	.clk(clk_clk),
	.d(\E_rot_step1[22]~18_combout ),
	.asdata(\E_rot_step1[26]~19_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add10~1_combout ),
	.ena(!\A_mem_stall~q ),
	.q(\M_rot_prestep2[26]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[26] .is_wysiwyg = "true";
defparam \M_rot_prestep2[26] .power_up = "low";

cyclonev_lcell_comb \M_rot[2]~16 (
	.dataa(!\M_rot_prestep2[10]~q ),
	.datab(!\M_rot_prestep2[2]~q ),
	.datac(!\M_rot_prestep2[26]~q ),
	.datad(!\M_rot_prestep2[18]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[2]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[2]~16 .extended_lut = "off";
defparam \M_rot[2]~16 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[2]~16 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~16 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_mask[2]~q ),
	.datac(!\M_rot_pass1~q ),
	.datad(!\M_rot_sel_fill1~q ),
	.datae(!\M_rot[2]~16_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~16 .extended_lut = "off";
defparam \A_shift_rot_result~16 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~16 .shared_arith = "off";

dffeas \A_shift_rot_result[10] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~16_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_shift_rot_result[10]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[10] .is_wysiwyg = "true";
defparam \A_shift_rot_result[10] .power_up = "low";

dffeas \A_inst_result[10] (
	.clk(clk_clk),
	.d(\M_pc_plus_one[8]~q ),
	.asdata(\M_alu_result[10]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\A_inst_result[9]~0_combout ),
	.sload(!\M_exc_any~combout ),
	.ena(!\A_mem_stall~q ),
	.q(\A_inst_result[10]~q ),
	.prn(vcc));
defparam \A_inst_result[10] .is_wysiwyg = "true";
defparam \A_inst_result[10] .power_up = "low";

dffeas \A_mul_cell_p1[10] (
	.clk(clk_clk),
	.d(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[10]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_mul_cell_p1[10]~q ),
	.prn(vcc));
defparam \A_mul_cell_p1[10] .is_wysiwyg = "true";
defparam \A_mul_cell_p1[10] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[10]~18 (
	.dataa(!\A_slow_inst_result[10]~q ),
	.datab(!\A_shift_rot_result[10]~q ),
	.datac(!\A_inst_result[10]~q ),
	.datad(!\A_mul_cell_p1[10]~q ),
	.datae(!\A_wr_data_unfiltered[15]~0_combout ),
	.dataf(!\A_wr_data_unfiltered[15]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[10]~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[10]~18 .extended_lut = "off";
defparam \A_wr_data_unfiltered[10]~18 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_wr_data_unfiltered[10]~18 .shared_arith = "off";

dffeas \W_wr_data[10] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[10]~18_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[10]~q ),
	.prn(vcc));
defparam \W_wr_data[10] .is_wysiwyg = "true";
defparam \W_wr_data[10] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[10]~43 (
	.dataa(!\D_src2_reg[0]~7_combout ),
	.datab(!\D_src2_reg[0]~8_combout ),
	.datac(!\W_wr_data[10]~q ),
	.datad(!\A_wr_data_unfiltered[10]~18_combout ),
	.datae(!\M_alu_result[10]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[10]~43_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[10]~43 .extended_lut = "off";
defparam \D_src2_reg[10]~43 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \D_src2_reg[10]~43 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[10]~44 (
	.dataa(!\D_src2_reg[0]~4_combout ),
	.datab(!\D_src2_reg[0]~5_combout ),
	.datac(!\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[10] ),
	.datad(!\E_alu_result[10]~combout ),
	.datae(!\D_src2_reg[10]~43_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[10]~44_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[10]~44 .extended_lut = "off";
defparam \D_src2_reg[10]~44 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \D_src2_reg[10]~44 .shared_arith = "off";

dffeas \E_src2[10] (
	.clk(clk_clk),
	.d(\D_iw[16]~q ),
	.asdata(\D_src2_reg[10]~44_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src2[5]~2_combout ),
	.sload(!\D_ctrl_src2_choose_imm~q ),
	.ena(!\A_mem_stall~q ),
	.q(\E_src2[10]~q ),
	.prn(vcc));
defparam \E_src2[10] .is_wysiwyg = "true";
defparam \E_src2[10] .power_up = "low";

cyclonev_lcell_comb \E_alu_result~13 (
	.dataa(!\E_src2[10]~q ),
	.datab(!\E_src1[10]~q ),
	.datac(!\E_logic_op[1]~q ),
	.datad(!\E_logic_op[0]~q ),
	.datae(!\E_ctrl_logic~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result~13 .extended_lut = "off";
defparam \E_alu_result~13 .lut_mask = 64'h6996FFFF6996FFFF;
defparam \E_alu_result~13 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[10] (
	.dataa(!\Add9~37_sumout ),
	.datab(!\E_ctrl_retaddr~q ),
	.datac(!\E_alu_result~0_combout ),
	.datad(!\E_alu_result~13_combout ),
	.datae(!\E_extra_pc[8]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[10]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[10] .extended_lut = "off";
defparam \E_alu_result[10] .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \E_alu_result[10] .shared_arith = "off";

dffeas \M_alu_result[10] (
	.clk(clk_clk),
	.d(\E_alu_result[10]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_alu_result[10]~q ),
	.prn(vcc));
defparam \M_alu_result[10] .is_wysiwyg = "true";
defparam \M_alu_result[10] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[10]~12 (
	.dataa(!\M_alu_result[10]~q ),
	.datab(!\A_wr_data_unfiltered[10]~18_combout ),
	.datac(!\first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[10] ),
	.datad(!\W_wr_data[10]~q ),
	.datae(!\E_src1[26]~0_combout ),
	.dataf(!\E_src1[26]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[10]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[10]~12 .extended_lut = "off";
defparam \D_src1_reg[10]~12 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[10]~12 .shared_arith = "off";

dffeas \E_src1[10] (
	.clk(clk_clk),
	.d(\D_src1_reg[10]~12_combout ),
	.asdata(\E_alu_result[10]~combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\Equal303~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(!\A_mem_stall~q ),
	.q(\E_src1[10]~q ),
	.prn(vcc));
defparam \E_src1[10] .is_wysiwyg = "true";
defparam \E_src1[10] .power_up = "low";

cyclonev_lcell_comb \E_rot_step1[10]~23 (
	.dataa(!\E_src1[10]~q ),
	.datab(!\E_src1[9]~q ),
	.datac(!\E_src1[8]~q ),
	.datad(!\E_src1[7]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add10~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[10]~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[10]~23 .extended_lut = "off";
defparam \E_rot_step1[10]~23 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[10]~23 .shared_arith = "off";

dffeas \M_rot_prestep2[14] (
	.clk(clk_clk),
	.d(\E_rot_step1[10]~23_combout ),
	.asdata(\E_rot_step1[14]~20_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add10~1_combout ),
	.ena(!\A_mem_stall~q ),
	.q(\M_rot_prestep2[14]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[14] .is_wysiwyg = "true";
defparam \M_rot_prestep2[14] .power_up = "low";

cyclonev_lcell_comb \M_rot[6]~30 (
	.dataa(!\M_rot_prestep2[14]~q ),
	.datab(!\M_rot_prestep2[6]~q ),
	.datac(!\M_rot_prestep2[30]~q ),
	.datad(!\M_rot_prestep2[22]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[6]~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[6]~30 .extended_lut = "off";
defparam \M_rot[6]~30 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[6]~30 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~30 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_mask[6]~q ),
	.datac(!\M_rot_pass1~q ),
	.datad(!\M_rot_sel_fill1~q ),
	.datae(!\M_rot[6]~30_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~30 .extended_lut = "off";
defparam \A_shift_rot_result~30 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~30 .shared_arith = "off";

dffeas \A_shift_rot_result[14] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~30_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_shift_rot_result[14]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[14] .is_wysiwyg = "true";
defparam \A_shift_rot_result[14] .power_up = "low";

dffeas \A_inst_result[14] (
	.clk(clk_clk),
	.d(\M_pc_plus_one[12]~q ),
	.asdata(\M_alu_result[14]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\A_inst_result[9]~0_combout ),
	.sload(!\M_exc_any~combout ),
	.ena(!\A_mem_stall~q ),
	.q(\A_inst_result[14]~q ),
	.prn(vcc));
defparam \A_inst_result[14] .is_wysiwyg = "true";
defparam \A_inst_result[14] .power_up = "low";

dffeas \A_mul_cell_p1[14] (
	.clk(clk_clk),
	.d(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[14]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_mul_cell_p1[14]~q ),
	.prn(vcc));
defparam \A_mul_cell_p1[14] .is_wysiwyg = "true";
defparam \A_mul_cell_p1[14] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[14]~32 (
	.dataa(!\A_slow_inst_result[14]~q ),
	.datab(!\A_shift_rot_result[14]~q ),
	.datac(!\A_inst_result[14]~q ),
	.datad(!\A_mul_cell_p1[14]~q ),
	.datae(!\A_wr_data_unfiltered[15]~0_combout ),
	.dataf(!\A_wr_data_unfiltered[15]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[14]~32_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[14]~32 .extended_lut = "off";
defparam \A_wr_data_unfiltered[14]~32 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_wr_data_unfiltered[14]~32 .shared_arith = "off";

dffeas \W_wr_data[14] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[14]~32_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[14]~q ),
	.prn(vcc));
defparam \W_wr_data[14] .is_wysiwyg = "true";
defparam \W_wr_data[14] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[14]~68 (
	.dataa(!\D_src2_reg[0]~7_combout ),
	.datab(!\D_src2_reg[0]~8_combout ),
	.datac(!\W_wr_data[14]~q ),
	.datad(!\A_wr_data_unfiltered[14]~32_combout ),
	.datae(!\M_alu_result[14]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[14]~68_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[14]~68 .extended_lut = "off";
defparam \D_src2_reg[14]~68 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \D_src2_reg[14]~68 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[14]~69 (
	.dataa(!\D_src2_reg[0]~4_combout ),
	.datab(!\D_src2_reg[0]~5_combout ),
	.datac(!\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[14] ),
	.datad(!\E_alu_result[14]~combout ),
	.datae(!\D_src2_reg[14]~68_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[14]~69_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[14]~69 .extended_lut = "off";
defparam \D_src2_reg[14]~69 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \D_src2_reg[14]~69 .shared_arith = "off";

dffeas \E_src2[14] (
	.clk(clk_clk),
	.d(\D_iw[20]~q ),
	.asdata(\D_src2_reg[14]~69_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src2[5]~2_combout ),
	.sload(!\D_ctrl_src2_choose_imm~q ),
	.ena(!\A_mem_stall~q ),
	.q(\E_src2[14]~q ),
	.prn(vcc));
defparam \E_src2[14] .is_wysiwyg = "true";
defparam \E_src2[14] .power_up = "low";

cyclonev_lcell_comb \E_alu_result~23 (
	.dataa(!\E_src2[14]~q ),
	.datab(!\E_src1[14]~q ),
	.datac(!\E_logic_op[1]~q ),
	.datad(!\E_logic_op[0]~q ),
	.datae(!\E_ctrl_logic~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result~23 .extended_lut = "off";
defparam \E_alu_result~23 .lut_mask = 64'h6996FFFF6996FFFF;
defparam \E_alu_result~23 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[14] (
	.dataa(!\Add9~21_sumout ),
	.datab(!\E_ctrl_retaddr~q ),
	.datac(!\E_alu_result~0_combout ),
	.datad(!\E_alu_result~23_combout ),
	.datae(!\E_extra_pc[12]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[14]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[14] .extended_lut = "off";
defparam \E_alu_result[14] .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \E_alu_result[14] .shared_arith = "off";

dffeas \M_alu_result[14] (
	.clk(clk_clk),
	.d(\E_alu_result[14]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_alu_result[14]~q ),
	.prn(vcc));
defparam \M_alu_result[14] .is_wysiwyg = "true";
defparam \M_alu_result[14] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[14]~30 (
	.dataa(!\M_alu_result[14]~q ),
	.datab(!\A_wr_data_unfiltered[14]~32_combout ),
	.datac(!\first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[14] ),
	.datad(!\W_wr_data[14]~q ),
	.datae(!\E_src1[26]~0_combout ),
	.dataf(!\E_src1[26]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[14]~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[14]~30 .extended_lut = "off";
defparam \D_src1_reg[14]~30 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[14]~30 .shared_arith = "off";

dffeas \E_src1[14] (
	.clk(clk_clk),
	.d(\D_src1_reg[14]~30_combout ),
	.asdata(\E_alu_result[14]~combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\Equal303~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(!\A_mem_stall~q ),
	.q(\E_src1[14]~q ),
	.prn(vcc));
defparam \E_src1[14] .is_wysiwyg = "true";
defparam \E_src1[14] .power_up = "low";

cyclonev_lcell_comb \E_rot_step1[14]~20 (
	.dataa(!\E_src1[14]~q ),
	.datab(!\E_src1[13]~q ),
	.datac(!\E_src1[12]~q ),
	.datad(!\E_src1[11]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add10~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[14]~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[14]~20 .extended_lut = "off";
defparam \E_rot_step1[14]~20 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[14]~20 .shared_arith = "off";

dffeas \M_rot_prestep2[18] (
	.clk(clk_clk),
	.d(\E_rot_step1[14]~20_combout ),
	.asdata(\E_rot_step1[18]~21_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add10~1_combout ),
	.ena(!\A_mem_stall~q ),
	.q(\M_rot_prestep2[18]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[18] .is_wysiwyg = "true";
defparam \M_rot_prestep2[18] .power_up = "low";

cyclonev_lcell_comb \M_rot[2]~25 (
	.dataa(!\M_rot_prestep2[18]~q ),
	.datab(!\M_rot_prestep2[10]~q ),
	.datac(!\M_rot_prestep2[2]~q ),
	.datad(!\M_rot_prestep2[26]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[2]~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[2]~25 .extended_lut = "off";
defparam \M_rot[2]~25 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[2]~25 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~25 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_mask[2]~q ),
	.datac(!\M_rot_pass2~q ),
	.datad(!\M_rot_sel_fill2~q ),
	.datae(!\M_rot[2]~25_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~25 .extended_lut = "off";
defparam \A_shift_rot_result~25 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~25 .shared_arith = "off";

dffeas \A_shift_rot_result[18] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~25_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_shift_rot_result[18]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[18] .is_wysiwyg = "true";
defparam \A_shift_rot_result[18] .power_up = "low";

dffeas \A_inst_result[18] (
	.clk(clk_clk),
	.d(\M_alu_result[18]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\A_inst_result[26]~1_combout ),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_inst_result[18]~q ),
	.prn(vcc));
defparam \A_inst_result[18] .is_wysiwyg = "true";
defparam \A_inst_result[18] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[18]~27 (
	.dataa(!\A_slow_inst_result[18]~q ),
	.datab(!\A_shift_rot_result[18]~q ),
	.datac(!\A_inst_result[18]~q ),
	.datad(!\Add12~53_sumout ),
	.datae(!\A_wr_data_unfiltered[15]~0_combout ),
	.dataf(!\A_wr_data_unfiltered[15]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[18]~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[18]~27 .extended_lut = "off";
defparam \A_wr_data_unfiltered[18]~27 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_wr_data_unfiltered[18]~27 .shared_arith = "off";

dffeas \W_wr_data[18] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[18]~27_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[18]~q ),
	.prn(vcc));
defparam \W_wr_data[18] .is_wysiwyg = "true";
defparam \W_wr_data[18] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[18]~60 (
	.dataa(!\D_src2_reg[0]~4_combout ),
	.datab(!\D_src2_reg[0]~7_combout ),
	.datac(!\D_src2_reg[0]~8_combout ),
	.datad(!\M_alu_result[18]~q ),
	.datae(!\A_wr_data_unfiltered[18]~27_combout ),
	.dataf(!\W_wr_data[18]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[18]~60_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[18]~60 .extended_lut = "off";
defparam \D_src2_reg[18]~60 .lut_mask = 64'hBEFFFFFFFFFFFFFF;
defparam \D_src2_reg[18]~60 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[18]~35 (
	.dataa(!\D_ctrl_hi_imm16~q ),
	.datab(!\D_iw[21]~q ),
	.datac(!\D_ctrl_unsigned_lo_imm16~q ),
	.datad(!\D_iw[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[18]~35_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[18]~35 .extended_lut = "off";
defparam \D_src2[18]~35 .lut_mask = 64'h7BFF7BFF7BFF7BFF;
defparam \D_src2[18]~35 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[18]~36 (
	.dataa(!\D_ctrl_src2_choose_imm~q ),
	.datab(!\E_logic_result[18]~11_combout ),
	.datac(!\E_ctrl_logic~q ),
	.datad(!\E_alu_result~0_combout ),
	.datae(!\Add9~125_sumout ),
	.dataf(!\D_src2[18]~35_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[18]~36_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[18]~36 .extended_lut = "off";
defparam \D_src2[18]~36 .lut_mask = 64'h27FFFFFFFFFFFFFF;
defparam \D_src2[18]~36 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[18]~25 (
	.dataa(!\D_src2_reg[0]~5_combout ),
	.datab(!\D_ctrl_src2_choose_imm~q ),
	.datac(!\D_src2_reg[18]~60_combout ),
	.datad(!\D_src2_reg[0]~4_combout ),
	.datae(!\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[18] ),
	.dataf(!\D_src2[18]~36_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[18]~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[18]~25 .extended_lut = "off";
defparam \D_src2[18]~25 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \D_src2[18]~25 .shared_arith = "off";

dffeas \E_src2[18] (
	.clk(clk_clk),
	.d(\D_src2[18]~25_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src2[30]~1_combout ),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_src2[18]~q ),
	.prn(vcc));
defparam \E_src2[18] .is_wysiwyg = "true";
defparam \E_src2[18] .power_up = "low";

cyclonev_lcell_comb \E_logic_result[18]~11 (
	.dataa(!\E_src2[18]~q ),
	.datab(!\E_src1[18]~q ),
	.datac(!\E_logic_op[1]~q ),
	.datad(!\E_logic_op[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[18]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[18]~11 .extended_lut = "off";
defparam \E_logic_result[18]~11 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[18]~11 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[18] (
	.dataa(!\E_logic_result[18]~11_combout ),
	.datab(!\E_ctrl_logic~q ),
	.datac(!\E_alu_result~0_combout ),
	.datad(!\Add9~125_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[18]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[18] .extended_lut = "off";
defparam \E_alu_result[18] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \E_alu_result[18] .shared_arith = "off";

dffeas \M_alu_result[18] (
	.clk(clk_clk),
	.d(\E_alu_result[18]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_alu_result[18]~q ),
	.prn(vcc));
defparam \M_alu_result[18] .is_wysiwyg = "true";
defparam \M_alu_result[18] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[18]~25 (
	.dataa(!\M_alu_result[18]~q ),
	.datab(!\A_wr_data_unfiltered[18]~27_combout ),
	.datac(!\first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[18] ),
	.datad(!\W_wr_data[18]~q ),
	.datae(!\E_src1[26]~0_combout ),
	.dataf(!\E_src1[26]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[18]~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[18]~25 .extended_lut = "off";
defparam \D_src1_reg[18]~25 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[18]~25 .shared_arith = "off";

dffeas \E_src1[18] (
	.clk(clk_clk),
	.d(\D_src1_reg[18]~25_combout ),
	.asdata(\E_alu_result[18]~combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\Equal303~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(!\A_mem_stall~q ),
	.q(\E_src1[18]~q ),
	.prn(vcc));
defparam \E_src1[18] .is_wysiwyg = "true";
defparam \E_src1[18] .power_up = "low";

cyclonev_lcell_comb \E_rot_step1[18]~21 (
	.dataa(!\E_src1[18]~q ),
	.datab(!\E_src1[17]~q ),
	.datac(!\E_src1[16]~q ),
	.datad(!\E_src1[15]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add10~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[18]~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[18]~21 .extended_lut = "off";
defparam \E_rot_step1[18]~21 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[18]~21 .shared_arith = "off";

dffeas \M_rot_prestep2[22] (
	.clk(clk_clk),
	.d(\E_rot_step1[18]~21_combout ),
	.asdata(\E_rot_step1[22]~18_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add10~1_combout ),
	.ena(!\A_mem_stall~q ),
	.q(\M_rot_prestep2[22]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[22] .is_wysiwyg = "true";
defparam \M_rot_prestep2[22] .power_up = "low";

cyclonev_lcell_comb \M_rot[6]~8 (
	.dataa(!\M_rot_prestep2[22]~q ),
	.datab(!\M_rot_prestep2[14]~q ),
	.datac(!\M_rot_prestep2[6]~q ),
	.datad(!\M_rot_prestep2[30]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[6]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[6]~8 .extended_lut = "off";
defparam \M_rot[6]~8 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[6]~8 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~8 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_mask[6]~q ),
	.datac(!\M_rot_pass2~q ),
	.datad(!\M_rot_sel_fill2~q ),
	.datae(!\M_rot[6]~8_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~8 .extended_lut = "off";
defparam \A_shift_rot_result~8 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~8 .shared_arith = "off";

dffeas \A_shift_rot_result[22] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~8_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_shift_rot_result[22]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[22] .is_wysiwyg = "true";
defparam \A_shift_rot_result[22] .power_up = "low";

dffeas \A_inst_result[22] (
	.clk(clk_clk),
	.d(\M_alu_result[22]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\A_inst_result[26]~1_combout ),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_inst_result[22]~q ),
	.prn(vcc));
defparam \A_inst_result[22] .is_wysiwyg = "true";
defparam \A_inst_result[22] .power_up = "low";

cyclonev_lcell_comb \Add11~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[6]~q ),
	.datae(gnd),
	.dataf(!\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[22]~q ),
	.datag(gnd),
	.cin(\Add11~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add11~1_sumout ),
	.cout(\Add11~2 ),
	.shareout());
defparam \Add11~1 .extended_lut = "off";
defparam \Add11~1 .lut_mask = 64'h0000FF00000000FF;
defparam \Add11~1 .shared_arith = "off";

dffeas \A_mul_s1[6] (
	.clk(clk_clk),
	.d(\Add11~1_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_mul_s1[6]~q ),
	.prn(vcc));
defparam \A_mul_s1[6] .is_wysiwyg = "true";
defparam \A_mul_s1[6] .power_up = "low";

dffeas \A_mul_cell_p3[6] (
	.clk(clk_clk),
	.d(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p3|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[6]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_mul_cell_p3[6]~q ),
	.prn(vcc));
defparam \A_mul_cell_p3[6] .is_wysiwyg = "true";
defparam \A_mul_cell_p3[6] .power_up = "low";

cyclonev_lcell_comb \Add12~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_mul_s1[6]~q ),
	.datae(gnd),
	.dataf(!\A_mul_cell_p3[6]~q ),
	.datag(gnd),
	.cin(\Add12~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add12~1_sumout ),
	.cout(\Add12~2 ),
	.shareout());
defparam \Add12~1 .extended_lut = "off";
defparam \Add12~1 .lut_mask = 64'h0000FF00000000FF;
defparam \Add12~1 .shared_arith = "off";

cyclonev_lcell_comb \A_wr_data_unfiltered[22]~10 (
	.dataa(!\A_slow_inst_result[22]~q ),
	.datab(!\A_shift_rot_result[22]~q ),
	.datac(!\A_inst_result[22]~q ),
	.datad(!\Add12~1_sumout ),
	.datae(!\A_wr_data_unfiltered[15]~0_combout ),
	.dataf(!\A_wr_data_unfiltered[15]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[22]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[22]~10 .extended_lut = "off";
defparam \A_wr_data_unfiltered[22]~10 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_wr_data_unfiltered[22]~10 .shared_arith = "off";

dffeas \W_wr_data[22] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[22]~10_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[22]~q ),
	.prn(vcc));
defparam \W_wr_data[22] .is_wysiwyg = "true";
defparam \W_wr_data[22] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[22]~1 (
	.dataa(!\M_alu_result[22]~q ),
	.datab(!\A_wr_data_unfiltered[22]~10_combout ),
	.datac(!\first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[22] ),
	.datad(!\W_wr_data[22]~q ),
	.datae(!\E_src1[26]~0_combout ),
	.dataf(!\E_src1[26]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[22]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[22]~1 .extended_lut = "off";
defparam \D_src1_reg[22]~1 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[22]~1 .shared_arith = "off";

dffeas \E_src1[22] (
	.clk(clk_clk),
	.d(\D_src1_reg[22]~1_combout ),
	.asdata(\E_alu_result[22]~combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\Equal303~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(!\A_mem_stall~q ),
	.q(\E_src1[22]~q ),
	.prn(vcc));
defparam \E_src1[22] .is_wysiwyg = "true";
defparam \E_src1[22] .power_up = "low";

cyclonev_lcell_comb \E_logic_result[22]~1 (
	.dataa(!\E_src2[22]~q ),
	.datab(!\E_src1[22]~q ),
	.datac(!\E_logic_op[1]~q ),
	.datad(!\E_logic_op[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[22]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[22]~1 .extended_lut = "off";
defparam \E_logic_result[22]~1 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[22]~1 .shared_arith = "off";

cyclonev_lcell_comb \Add9~77 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[22]~q ),
	.datae(gnd),
	.dataf(!\E_src1[22]~q ),
	.datag(gnd),
	.cin(\Add9~94 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~77_sumout ),
	.cout(\Add9~78 ),
	.shareout());
defparam \Add9~77 .extended_lut = "off";
defparam \Add9~77 .lut_mask = 64'h0000FF00000055AA;
defparam \Add9~77 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[22] (
	.dataa(!\E_logic_result[22]~1_combout ),
	.datab(!\E_ctrl_logic~q ),
	.datac(!\E_alu_result~0_combout ),
	.datad(!\Add9~77_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[22]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[22] .extended_lut = "off";
defparam \E_alu_result[22] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \E_alu_result[22] .shared_arith = "off";

dffeas \M_alu_result[22] (
	.clk(clk_clk),
	.d(\E_alu_result[22]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_alu_result[22]~q ),
	.prn(vcc));
defparam \M_alu_result[22] .is_wysiwyg = "true";
defparam \M_alu_result[22] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[22]~26 (
	.dataa(!\D_src2_reg[0]~4_combout ),
	.datab(!\D_src2_reg[0]~7_combout ),
	.datac(!\D_src2_reg[0]~8_combout ),
	.datad(!\M_alu_result[22]~q ),
	.datae(!\A_wr_data_unfiltered[22]~10_combout ),
	.dataf(!\W_wr_data[22]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[22]~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[22]~26 .extended_lut = "off";
defparam \D_src2_reg[22]~26 .lut_mask = 64'hBEFFFFFFFFFFFFFF;
defparam \D_src2_reg[22]~26 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[22]~41 (
	.dataa(!\D_iw[12]~q ),
	.datab(!\D_ctrl_hi_imm16~q ),
	.datac(!\D_iw[21]~q ),
	.datad(!\D_ctrl_unsigned_lo_imm16~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[22]~41_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[22]~41 .extended_lut = "off";
defparam \D_src2[22]~41 .lut_mask = 64'h7FDF7FDF7FDF7FDF;
defparam \D_src2[22]~41 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[22]~42 (
	.dataa(!\D_ctrl_src2_choose_imm~q ),
	.datab(!\E_logic_result[22]~1_combout ),
	.datac(!\E_ctrl_logic~q ),
	.datad(!\E_alu_result~0_combout ),
	.datae(!\Add9~77_sumout ),
	.dataf(!\D_src2[22]~41_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[22]~42_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[22]~42 .extended_lut = "off";
defparam \D_src2[22]~42 .lut_mask = 64'h27FFFFFFFFFFFFFF;
defparam \D_src2[22]~42 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[22]~1 (
	.dataa(!\D_src2_reg[0]~5_combout ),
	.datab(!\D_ctrl_src2_choose_imm~q ),
	.datac(!\D_src2_reg[22]~26_combout ),
	.datad(!\D_src2_reg[0]~4_combout ),
	.datae(!\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[22] ),
	.dataf(!\D_src2[22]~42_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[22]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[22]~1 .extended_lut = "off";
defparam \D_src2[22]~1 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \D_src2[22]~1 .shared_arith = "off";

dffeas \E_src2[22] (
	.clk(clk_clk),
	.d(\D_src2[22]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src2[30]~1_combout ),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_src2[22]~q ),
	.prn(vcc));
defparam \E_src2[22] .is_wysiwyg = "true";
defparam \E_src2[22] .power_up = "low";

cyclonev_lcell_comb \Add9~81 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[23]~q ),
	.datae(gnd),
	.dataf(!\E_src1[23]~q ),
	.datag(gnd),
	.cin(\Add9~78 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~81_sumout ),
	.cout(\Add9~82 ),
	.shareout());
defparam \Add9~81 .extended_lut = "off";
defparam \Add9~81 .lut_mask = 64'h0000FF00000055AA;
defparam \Add9~81 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[23] (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\E_alu_result~7_combout ),
	.datac(!\Add9~81_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[23]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[23] .extended_lut = "off";
defparam \E_alu_result[23] .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \E_alu_result[23] .shared_arith = "off";

dffeas \M_alu_result[23] (
	.clk(clk_clk),
	.d(\E_alu_result[23]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_alu_result[23]~q ),
	.prn(vcc));
defparam \M_alu_result[23] .is_wysiwyg = "true";
defparam \M_alu_result[23] .power_up = "low";

cyclonev_lcell_comb \A_slow_inst_result_nxt[23]~36 (
	.dataa(!\A_ctrl_ld32~q ),
	.datab(!\A_ld_align_byte2_byte3_fill~q ),
	.datac(!src0_valid),
	.datad(!av_readdata_pre_23),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[23]~36_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[23]~36 .extended_lut = "off";
defparam \A_slow_inst_result_nxt[23]~36 .lut_mask = 64'h27FF27FF27FF27FF;
defparam \A_slow_inst_result_nxt[23]~36 .shared_arith = "off";

cyclonev_lcell_comb \A_slow_inst_result_nxt[23]~9 (
	.dataa(!\A_ctrl_ld32~q ),
	.datab(!\d_readdata_d1[23]~q ),
	.datac(!\A_slow_ld_data_fill_bit~0_combout ),
	.datad(!src0_valid1),
	.datae(!q_a_23),
	.dataf(!\A_slow_inst_result_nxt[23]~36_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[23]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[23]~9 .extended_lut = "off";
defparam \A_slow_inst_result_nxt[23]~9 .lut_mask = 64'h7FFFFFFFBFFFFFFF;
defparam \A_slow_inst_result_nxt[23]~9 .shared_arith = "off";

dffeas \A_slow_inst_result[23] (
	.clk(clk_clk),
	.d(\A_slow_inst_result_nxt[23]~9_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_ctrl_ld~q ),
	.q(\A_slow_inst_result[23]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[23] .is_wysiwyg = "true";
defparam \A_slow_inst_result[23] .power_up = "low";

cyclonev_lcell_comb \M_rot[7]~9 (
	.dataa(!\M_rot_prestep2[23]~q ),
	.datab(!\M_rot_prestep2[15]~q ),
	.datac(!\M_rot_prestep2[7]~q ),
	.datad(!\M_rot_prestep2[31]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[7]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[7]~9 .extended_lut = "off";
defparam \M_rot[7]~9 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[7]~9 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~9 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_mask[7]~q ),
	.datac(!\M_rot_pass2~q ),
	.datad(!\M_rot_sel_fill2~q ),
	.datae(!\M_rot[7]~9_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~9 .extended_lut = "off";
defparam \A_shift_rot_result~9 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~9 .shared_arith = "off";

dffeas \A_shift_rot_result[23] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~9_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_shift_rot_result[23]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[23] .is_wysiwyg = "true";
defparam \A_shift_rot_result[23] .power_up = "low";

dffeas \A_inst_result[23] (
	.clk(clk_clk),
	.d(\M_alu_result[23]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\A_inst_result[26]~1_combout ),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_inst_result[23]~q ),
	.prn(vcc));
defparam \A_inst_result[23] .is_wysiwyg = "true";
defparam \A_inst_result[23] .power_up = "low";

cyclonev_lcell_comb \Add11~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[7]~q ),
	.datae(gnd),
	.dataf(!\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[23]~q ),
	.datag(gnd),
	.cin(\Add11~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add11~5_sumout ),
	.cout(\Add11~6 ),
	.shareout());
defparam \Add11~5 .extended_lut = "off";
defparam \Add11~5 .lut_mask = 64'h0000FF00000000FF;
defparam \Add11~5 .shared_arith = "off";

dffeas \A_mul_s1[7] (
	.clk(clk_clk),
	.d(\Add11~5_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_mul_s1[7]~q ),
	.prn(vcc));
defparam \A_mul_s1[7] .is_wysiwyg = "true";
defparam \A_mul_s1[7] .power_up = "low";

dffeas \A_mul_cell_p3[7] (
	.clk(clk_clk),
	.d(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p3|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[7]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_mul_cell_p3[7]~q ),
	.prn(vcc));
defparam \A_mul_cell_p3[7] .is_wysiwyg = "true";
defparam \A_mul_cell_p3[7] .power_up = "low";

cyclonev_lcell_comb \Add12~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_mul_s1[7]~q ),
	.datae(gnd),
	.dataf(!\A_mul_cell_p3[7]~q ),
	.datag(gnd),
	.cin(\Add12~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add12~5_sumout ),
	.cout(\Add12~6 ),
	.shareout());
defparam \Add12~5 .extended_lut = "off";
defparam \Add12~5 .lut_mask = 64'h0000FF00000000FF;
defparam \Add12~5 .shared_arith = "off";

cyclonev_lcell_comb \A_wr_data_unfiltered[23]~11 (
	.dataa(!\A_slow_inst_result[23]~q ),
	.datab(!\A_shift_rot_result[23]~q ),
	.datac(!\A_inst_result[23]~q ),
	.datad(!\Add12~5_sumout ),
	.datae(!\A_wr_data_unfiltered[15]~0_combout ),
	.dataf(!\A_wr_data_unfiltered[15]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[23]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[23]~11 .extended_lut = "off";
defparam \A_wr_data_unfiltered[23]~11 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_wr_data_unfiltered[23]~11 .shared_arith = "off";

dffeas \W_wr_data[23] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[23]~11_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[23]~q ),
	.prn(vcc));
defparam \W_wr_data[23] .is_wysiwyg = "true";
defparam \W_wr_data[23] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[23]~2 (
	.dataa(!\M_alu_result[23]~q ),
	.datab(!\A_wr_data_unfiltered[23]~11_combout ),
	.datac(!\first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[23] ),
	.datad(!\W_wr_data[23]~q ),
	.datae(!\E_src1[26]~0_combout ),
	.dataf(!\E_src1[26]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[23]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[23]~2 .extended_lut = "off";
defparam \D_src1_reg[23]~2 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[23]~2 .shared_arith = "off";

dffeas \E_src1[23] (
	.clk(clk_clk),
	.d(\D_src1_reg[23]~2_combout ),
	.asdata(\E_alu_result[23]~combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\Equal303~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(!\A_mem_stall~q ),
	.q(\E_src1[23]~q ),
	.prn(vcc));
defparam \E_src1[23] .is_wysiwyg = "true";
defparam \E_src1[23] .power_up = "low";

cyclonev_lcell_comb \E_logic_result[23]~2 (
	.dataa(!\E_src2[23]~q ),
	.datab(!\E_src1[23]~q ),
	.datac(!\E_logic_op[1]~q ),
	.datad(!\E_logic_op[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[23]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[23]~2 .extended_lut = "off";
defparam \E_logic_result[23]~2 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[23]~2 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result~7 (
	.dataa(!\E_logic_result[23]~2_combout ),
	.datab(!\E_ctrl_logic~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result~7 .extended_lut = "off";
defparam \E_alu_result~7 .lut_mask = 64'h7777777777777777;
defparam \E_alu_result~7 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[23]~27 (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\D_src2_reg[0]~2_combout ),
	.datac(!\E_alu_result~7_combout ),
	.datad(!\Add9~81_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[23]~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[23]~27 .extended_lut = "off";
defparam \D_src2_reg[23]~27 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \D_src2_reg[23]~27 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[0]~9 (
	.dataa(!\Equal304~0_combout ),
	.datab(!\D_src2_reg[0]~0_combout ),
	.datac(!\D_src2_reg[0]~1_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[0]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[0]~9 .extended_lut = "off";
defparam \D_src2_reg[0]~9 .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \D_src2_reg[0]~9 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[23]~28 (
	.dataa(!\D_src2_reg[0]~7_combout ),
	.datab(!\D_src2_reg[0]~8_combout ),
	.datac(!\D_src2_reg[0]~9_combout ),
	.datad(!\M_alu_result[23]~q ),
	.datae(!\A_wr_data_unfiltered[23]~11_combout ),
	.dataf(!\W_wr_data[23]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[23]~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[23]~28 .extended_lut = "off";
defparam \D_src2_reg[23]~28 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \D_src2_reg[23]~28 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[23]~2 (
	.dataa(!\D_iw[13]~q ),
	.datab(!\D_ctrl_hi_imm16~q ),
	.datac(!\D_iw[21]~q ),
	.datad(!\D_ctrl_unsigned_lo_imm16~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[23]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[23]~2 .extended_lut = "off";
defparam \D_src2[23]~2 .lut_mask = 64'h7FDF7FDF7FDF7FDF;
defparam \D_src2[23]~2 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[23]~3 (
	.dataa(!\D_src2_reg[0]~6_combout ),
	.datab(!\D_ctrl_src2_choose_imm~q ),
	.datac(!\D_src2_reg[23]~27_combout ),
	.datad(!\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[23] ),
	.datae(!\D_src2_reg[23]~28_combout ),
	.dataf(!\D_src2[23]~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[23]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[23]~3 .extended_lut = "off";
defparam \D_src2[23]~3 .lut_mask = 64'h47FFFFFFFFFFFFFF;
defparam \D_src2[23]~3 .shared_arith = "off";

dffeas \E_src2[23] (
	.clk(clk_clk),
	.d(\D_src2[23]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src2[30]~1_combout ),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_src2[23]~q ),
	.prn(vcc));
defparam \E_src2[23] .is_wysiwyg = "true";
defparam \E_src2[23] .power_up = "low";

cyclonev_lcell_comb \Add9~85 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[24]~q ),
	.datae(gnd),
	.dataf(!\E_src1[24]~q ),
	.datag(gnd),
	.cin(\Add9~82 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~85_sumout ),
	.cout(\Add9~86 ),
	.shareout());
defparam \Add9~85 .extended_lut = "off";
defparam \Add9~85 .lut_mask = 64'h0000FF00000055AA;
defparam \Add9~85 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[24] (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\E_alu_result~8_combout ),
	.datac(!\Add9~85_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[24]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[24] .extended_lut = "off";
defparam \E_alu_result[24] .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \E_alu_result[24] .shared_arith = "off";

dffeas \M_alu_result[24] (
	.clk(clk_clk),
	.d(\E_alu_result[24]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_alu_result[24]~q ),
	.prn(vcc));
defparam \M_alu_result[24] .is_wysiwyg = "true";
defparam \M_alu_result[24] .power_up = "low";

cyclonev_lcell_comb \A_slow_inst_result_nxt[24]~37 (
	.dataa(!\A_ctrl_ld32~q ),
	.datab(!\A_ld_align_byte2_byte3_fill~q ),
	.datac(!src0_valid),
	.datad(!av_readdata_pre_24),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[24]~37_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[24]~37 .extended_lut = "off";
defparam \A_slow_inst_result_nxt[24]~37 .lut_mask = 64'h27FF27FF27FF27FF;
defparam \A_slow_inst_result_nxt[24]~37 .shared_arith = "off";

cyclonev_lcell_comb \A_slow_inst_result_nxt[24]~10 (
	.dataa(!\A_ctrl_ld32~q ),
	.datab(!\d_readdata_d1[24]~q ),
	.datac(!\A_slow_ld_data_fill_bit~0_combout ),
	.datad(!src0_valid1),
	.datae(!q_a_24),
	.dataf(!\A_slow_inst_result_nxt[24]~37_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[24]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[24]~10 .extended_lut = "off";
defparam \A_slow_inst_result_nxt[24]~10 .lut_mask = 64'h7FFFFFFFBFFFFFFF;
defparam \A_slow_inst_result_nxt[24]~10 .shared_arith = "off";

dffeas \A_slow_inst_result[24] (
	.clk(clk_clk),
	.d(\A_slow_inst_result_nxt[24]~10_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_ctrl_ld~q ),
	.q(\A_slow_inst_result[24]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[24] .is_wysiwyg = "true";
defparam \A_slow_inst_result[24] .power_up = "low";

cyclonev_lcell_comb \E_rot_pass3~0 (
	.dataa(!\E_src2[3]~q ),
	.datab(!\E_src2[4]~q ),
	.datac(!\E_ctrl_rot~q ),
	.datad(!\E_ctrl_shift_rot_left~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_pass3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_pass3~0 .extended_lut = "off";
defparam \E_rot_pass3~0 .lut_mask = 64'hEFFFEFFFEFFFEFFF;
defparam \E_rot_pass3~0 .shared_arith = "off";

dffeas M_rot_pass3(
	.clk(clk_clk),
	.d(\E_rot_pass3~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_rot_pass3~q ),
	.prn(vcc));
defparam M_rot_pass3.is_wysiwyg = "true";
defparam M_rot_pass3.power_up = "low";

cyclonev_lcell_comb \E_rot_sel_fill3~0 (
	.dataa(!\E_src2[3]~q ),
	.datab(!\E_src2[4]~q ),
	.datac(!\E_ctrl_shift_rot_right~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_sel_fill3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_sel_fill3~0 .extended_lut = "off";
defparam \E_rot_sel_fill3~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \E_rot_sel_fill3~0 .shared_arith = "off";

dffeas M_rot_sel_fill3(
	.clk(clk_clk),
	.d(\E_rot_sel_fill3~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_rot_sel_fill3~q ),
	.prn(vcc));
defparam M_rot_sel_fill3.is_wysiwyg = "true";
defparam M_rot_sel_fill3.power_up = "low";

cyclonev_lcell_comb \M_rot[0]~10 (
	.dataa(!\M_rot_prestep2[24]~q ),
	.datab(!\M_rot_prestep2[16]~q ),
	.datac(!\M_rot_prestep2[8]~q ),
	.datad(!\M_rot_prestep2[0]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[0]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[0]~10 .extended_lut = "off";
defparam \M_rot[0]~10 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[0]~10 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~10 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_mask[0]~q ),
	.datac(!\M_rot_pass3~q ),
	.datad(!\M_rot_sel_fill3~q ),
	.datae(!\M_rot[0]~10_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~10 .extended_lut = "off";
defparam \A_shift_rot_result~10 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~10 .shared_arith = "off";

dffeas \A_shift_rot_result[24] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~10_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_shift_rot_result[24]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[24] .is_wysiwyg = "true";
defparam \A_shift_rot_result[24] .power_up = "low";

dffeas \A_inst_result[24] (
	.clk(clk_clk),
	.d(\M_alu_result[24]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\A_inst_result[26]~1_combout ),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_inst_result[24]~q ),
	.prn(vcc));
defparam \A_inst_result[24] .is_wysiwyg = "true";
defparam \A_inst_result[24] .power_up = "low";

cyclonev_lcell_comb \Add11~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[8]~q ),
	.datae(gnd),
	.dataf(!\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[24]~q ),
	.datag(gnd),
	.cin(\Add11~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add11~9_sumout ),
	.cout(\Add11~10 ),
	.shareout());
defparam \Add11~9 .extended_lut = "off";
defparam \Add11~9 .lut_mask = 64'h0000FF00000000FF;
defparam \Add11~9 .shared_arith = "off";

dffeas \A_mul_s1[8] (
	.clk(clk_clk),
	.d(\Add11~9_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_mul_s1[8]~q ),
	.prn(vcc));
defparam \A_mul_s1[8] .is_wysiwyg = "true";
defparam \A_mul_s1[8] .power_up = "low";

dffeas \A_mul_cell_p3[8] (
	.clk(clk_clk),
	.d(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p3|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[8]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_mul_cell_p3[8]~q ),
	.prn(vcc));
defparam \A_mul_cell_p3[8] .is_wysiwyg = "true";
defparam \A_mul_cell_p3[8] .power_up = "low";

cyclonev_lcell_comb \Add12~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_mul_s1[8]~q ),
	.datae(gnd),
	.dataf(!\A_mul_cell_p3[8]~q ),
	.datag(gnd),
	.cin(\Add12~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add12~9_sumout ),
	.cout(\Add12~10 ),
	.shareout());
defparam \Add12~9 .extended_lut = "off";
defparam \Add12~9 .lut_mask = 64'h0000FF00000000FF;
defparam \Add12~9 .shared_arith = "off";

cyclonev_lcell_comb \A_wr_data_unfiltered[24]~12 (
	.dataa(!\A_slow_inst_result[24]~q ),
	.datab(!\A_shift_rot_result[24]~q ),
	.datac(!\A_inst_result[24]~q ),
	.datad(!\Add12~9_sumout ),
	.datae(!\A_wr_data_unfiltered[15]~0_combout ),
	.dataf(!\A_wr_data_unfiltered[15]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[24]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[24]~12 .extended_lut = "off";
defparam \A_wr_data_unfiltered[24]~12 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_wr_data_unfiltered[24]~12 .shared_arith = "off";

dffeas \W_wr_data[24] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[24]~12_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[24]~q ),
	.prn(vcc));
defparam \W_wr_data[24] .is_wysiwyg = "true";
defparam \W_wr_data[24] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[24]~3 (
	.dataa(!\M_alu_result[24]~q ),
	.datab(!\A_wr_data_unfiltered[24]~12_combout ),
	.datac(!\first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[24] ),
	.datad(!\W_wr_data[24]~q ),
	.datae(!\E_src1[26]~0_combout ),
	.dataf(!\E_src1[26]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[24]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[24]~3 .extended_lut = "off";
defparam \D_src1_reg[24]~3 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[24]~3 .shared_arith = "off";

dffeas \E_src1[24] (
	.clk(clk_clk),
	.d(\D_src1_reg[24]~3_combout ),
	.asdata(\E_alu_result[24]~combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\Equal303~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(!\A_mem_stall~q ),
	.q(\E_src1[24]~q ),
	.prn(vcc));
defparam \E_src1[24] .is_wysiwyg = "true";
defparam \E_src1[24] .power_up = "low";

cyclonev_lcell_comb \E_logic_result[24]~3 (
	.dataa(!\E_src2[24]~q ),
	.datab(!\E_src1[24]~q ),
	.datac(!\E_logic_op[1]~q ),
	.datad(!\E_logic_op[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[24]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[24]~3 .extended_lut = "off";
defparam \E_logic_result[24]~3 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[24]~3 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result~8 (
	.dataa(!\E_logic_result[24]~3_combout ),
	.datab(!\E_ctrl_logic~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result~8 .extended_lut = "off";
defparam \E_alu_result~8 .lut_mask = 64'h7777777777777777;
defparam \E_alu_result~8 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[24]~29 (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\D_src2_reg[0]~2_combout ),
	.datac(!\E_alu_result~8_combout ),
	.datad(!\Add9~85_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[24]~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[24]~29 .extended_lut = "off";
defparam \D_src2_reg[24]~29 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \D_src2_reg[24]~29 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[24]~30 (
	.dataa(!\D_src2_reg[0]~7_combout ),
	.datab(!\D_src2_reg[0]~8_combout ),
	.datac(!\D_src2_reg[0]~9_combout ),
	.datad(!\M_alu_result[24]~q ),
	.datae(!\A_wr_data_unfiltered[24]~12_combout ),
	.dataf(!\W_wr_data[24]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[24]~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[24]~30 .extended_lut = "off";
defparam \D_src2_reg[24]~30 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \D_src2_reg[24]~30 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[24]~4 (
	.dataa(!\D_iw[14]~q ),
	.datab(!\D_ctrl_hi_imm16~q ),
	.datac(!\D_iw[21]~q ),
	.datad(!\D_ctrl_unsigned_lo_imm16~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[24]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[24]~4 .extended_lut = "off";
defparam \D_src2[24]~4 .lut_mask = 64'h7FDF7FDF7FDF7FDF;
defparam \D_src2[24]~4 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[24]~5 (
	.dataa(!\D_src2_reg[0]~6_combout ),
	.datab(!\D_ctrl_src2_choose_imm~q ),
	.datac(!\D_src2_reg[24]~29_combout ),
	.datad(!\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[24] ),
	.datae(!\D_src2_reg[24]~30_combout ),
	.dataf(!\D_src2[24]~4_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[24]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[24]~5 .extended_lut = "off";
defparam \D_src2[24]~5 .lut_mask = 64'h47FFFFFFFFFFFFFF;
defparam \D_src2[24]~5 .shared_arith = "off";

dffeas \E_src2[24] (
	.clk(clk_clk),
	.d(\D_src2[24]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src2[30]~1_combout ),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_src2[24]~q ),
	.prn(vcc));
defparam \E_src2[24] .is_wysiwyg = "true";
defparam \E_src2[24] .power_up = "low";

cyclonev_lcell_comb \Add9~89 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[25]~q ),
	.datae(gnd),
	.dataf(!\E_src1[25]~q ),
	.datag(gnd),
	.cin(\Add9~86 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~89_sumout ),
	.cout(\Add9~90 ),
	.shareout());
defparam \Add9~89 .extended_lut = "off";
defparam \Add9~89 .lut_mask = 64'h0000FF00000055AA;
defparam \Add9~89 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[25] (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\E_alu_result~9_combout ),
	.datac(!\Add9~89_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[25]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[25] .extended_lut = "off";
defparam \E_alu_result[25] .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \E_alu_result[25] .shared_arith = "off";

dffeas \M_alu_result[25] (
	.clk(clk_clk),
	.d(\E_alu_result[25]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_alu_result[25]~q ),
	.prn(vcc));
defparam \M_alu_result[25] .is_wysiwyg = "true";
defparam \M_alu_result[25] .power_up = "low";

cyclonev_lcell_comb \A_slow_inst_result_nxt[25]~39 (
	.dataa(!\A_ctrl_ld32~q ),
	.datab(!\A_ld_align_byte2_byte3_fill~q ),
	.datac(!src0_valid),
	.datad(!src_payload2),
	.datae(!av_readdata_pre_25),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[25]~39_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[25]~39 .extended_lut = "off";
defparam \A_slow_inst_result_nxt[25]~39 .lut_mask = 64'hFFFFFFD8FFFFFFD8;
defparam \A_slow_inst_result_nxt[25]~39 .shared_arith = "off";

cyclonev_lcell_comb \A_slow_inst_result_nxt[25]~11 (
	.dataa(!\A_ctrl_ld32~q ),
	.datab(!\d_readdata_d1[25]~q ),
	.datac(!\A_slow_ld_data_fill_bit~0_combout ),
	.datad(!src0_valid1),
	.datae(!q_a_25),
	.dataf(!\A_slow_inst_result_nxt[25]~39_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[25]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[25]~11 .extended_lut = "off";
defparam \A_slow_inst_result_nxt[25]~11 .lut_mask = 64'h7FFFFFFFBFFFFFFF;
defparam \A_slow_inst_result_nxt[25]~11 .shared_arith = "off";

dffeas \A_slow_inst_result[25] (
	.clk(clk_clk),
	.d(\A_slow_inst_result_nxt[25]~11_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_ctrl_ld~q ),
	.q(\A_slow_inst_result[25]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[25] .is_wysiwyg = "true";
defparam \A_slow_inst_result[25] .power_up = "low";

cyclonev_lcell_comb \M_rot[1]~11 (
	.dataa(!\M_rot_prestep2[25]~q ),
	.datab(!\M_rot_prestep2[17]~q ),
	.datac(!\M_rot_prestep2[9]~q ),
	.datad(!\M_rot_prestep2[1]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[1]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[1]~11 .extended_lut = "off";
defparam \M_rot[1]~11 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[1]~11 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~11 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_mask[1]~q ),
	.datac(!\M_rot_pass3~q ),
	.datad(!\M_rot_sel_fill3~q ),
	.datae(!\M_rot[1]~11_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~11 .extended_lut = "off";
defparam \A_shift_rot_result~11 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~11 .shared_arith = "off";

dffeas \A_shift_rot_result[25] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~11_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_shift_rot_result[25]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[25] .is_wysiwyg = "true";
defparam \A_shift_rot_result[25] .power_up = "low";

dffeas \A_inst_result[25] (
	.clk(clk_clk),
	.d(\M_alu_result[25]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\A_inst_result[26]~1_combout ),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_inst_result[25]~q ),
	.prn(vcc));
defparam \A_inst_result[25] .is_wysiwyg = "true";
defparam \A_inst_result[25] .power_up = "low";

cyclonev_lcell_comb \Add11~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[9]~q ),
	.datae(gnd),
	.dataf(!\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[25]~q ),
	.datag(gnd),
	.cin(\Add11~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add11~13_sumout ),
	.cout(\Add11~14 ),
	.shareout());
defparam \Add11~13 .extended_lut = "off";
defparam \Add11~13 .lut_mask = 64'h0000FF00000000FF;
defparam \Add11~13 .shared_arith = "off";

dffeas \A_mul_s1[9] (
	.clk(clk_clk),
	.d(\Add11~13_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_mul_s1[9]~q ),
	.prn(vcc));
defparam \A_mul_s1[9] .is_wysiwyg = "true";
defparam \A_mul_s1[9] .power_up = "low";

dffeas \A_mul_cell_p3[9] (
	.clk(clk_clk),
	.d(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p3|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[9]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_mul_cell_p3[9]~q ),
	.prn(vcc));
defparam \A_mul_cell_p3[9] .is_wysiwyg = "true";
defparam \A_mul_cell_p3[9] .power_up = "low";

cyclonev_lcell_comb \Add12~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_mul_s1[9]~q ),
	.datae(gnd),
	.dataf(!\A_mul_cell_p3[9]~q ),
	.datag(gnd),
	.cin(\Add12~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add12~13_sumout ),
	.cout(\Add12~14 ),
	.shareout());
defparam \Add12~13 .extended_lut = "off";
defparam \Add12~13 .lut_mask = 64'h0000FF00000000FF;
defparam \Add12~13 .shared_arith = "off";

cyclonev_lcell_comb \A_wr_data_unfiltered[25]~13 (
	.dataa(!\A_slow_inst_result[25]~q ),
	.datab(!\A_shift_rot_result[25]~q ),
	.datac(!\A_inst_result[25]~q ),
	.datad(!\Add12~13_sumout ),
	.datae(!\A_wr_data_unfiltered[15]~0_combout ),
	.dataf(!\A_wr_data_unfiltered[15]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[25]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[25]~13 .extended_lut = "off";
defparam \A_wr_data_unfiltered[25]~13 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_wr_data_unfiltered[25]~13 .shared_arith = "off";

dffeas \W_wr_data[25] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[25]~13_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[25]~q ),
	.prn(vcc));
defparam \W_wr_data[25] .is_wysiwyg = "true";
defparam \W_wr_data[25] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[25]~5 (
	.dataa(!\M_alu_result[25]~q ),
	.datab(!\A_wr_data_unfiltered[25]~13_combout ),
	.datac(!\first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[25] ),
	.datad(!\W_wr_data[25]~q ),
	.datae(!\E_src1[26]~0_combout ),
	.dataf(!\E_src1[26]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[25]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[25]~5 .extended_lut = "off";
defparam \D_src1_reg[25]~5 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[25]~5 .shared_arith = "off";

dffeas \E_src1[25] (
	.clk(clk_clk),
	.d(\D_src1_reg[25]~5_combout ),
	.asdata(\E_alu_result[25]~combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\Equal303~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(!\A_mem_stall~q ),
	.q(\E_src1[25]~q ),
	.prn(vcc));
defparam \E_src1[25] .is_wysiwyg = "true";
defparam \E_src1[25] .power_up = "low";

cyclonev_lcell_comb \E_alu_result~9 (
	.dataa(!\E_src2[25]~q ),
	.datab(!\E_src1[25]~q ),
	.datac(!\E_logic_op[1]~q ),
	.datad(!\E_logic_op[0]~q ),
	.datae(!\E_ctrl_logic~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result~9 .extended_lut = "off";
defparam \E_alu_result~9 .lut_mask = 64'h6996FFFF6996FFFF;
defparam \E_alu_result~9 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[25]~31 (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\D_src2_reg[0]~2_combout ),
	.datac(!\E_alu_result~9_combout ),
	.datad(!\Add9~89_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[25]~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[25]~31 .extended_lut = "off";
defparam \D_src2_reg[25]~31 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \D_src2_reg[25]~31 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[25]~32 (
	.dataa(!\D_src2_reg[0]~7_combout ),
	.datab(!\D_src2_reg[0]~8_combout ),
	.datac(!\D_src2_reg[0]~9_combout ),
	.datad(!\M_alu_result[25]~q ),
	.datae(!\A_wr_data_unfiltered[25]~13_combout ),
	.dataf(!\W_wr_data[25]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[25]~32_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[25]~32 .extended_lut = "off";
defparam \D_src2_reg[25]~32 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \D_src2_reg[25]~32 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[25]~6 (
	.dataa(!\D_iw[15]~q ),
	.datab(!\D_ctrl_hi_imm16~q ),
	.datac(!\D_iw[21]~q ),
	.datad(!\D_ctrl_unsigned_lo_imm16~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[25]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[25]~6 .extended_lut = "off";
defparam \D_src2[25]~6 .lut_mask = 64'h7FDF7FDF7FDF7FDF;
defparam \D_src2[25]~6 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[25]~7 (
	.dataa(!\D_src2_reg[0]~6_combout ),
	.datab(!\D_ctrl_src2_choose_imm~q ),
	.datac(!\D_src2_reg[25]~31_combout ),
	.datad(!\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[25] ),
	.datae(!\D_src2_reg[25]~32_combout ),
	.dataf(!\D_src2[25]~6_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[25]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[25]~7 .extended_lut = "off";
defparam \D_src2[25]~7 .lut_mask = 64'h47FFFFFFFFFFFFFF;
defparam \D_src2[25]~7 .shared_arith = "off";

dffeas \E_src2[25] (
	.clk(clk_clk),
	.d(\D_src2[25]~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src2[30]~1_combout ),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_src2[25]~q ),
	.prn(vcc));
defparam \E_src2[25] .is_wysiwyg = "true";
defparam \E_src2[25] .power_up = "low";

cyclonev_lcell_comb \Add9~105 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[26]~q ),
	.datae(gnd),
	.dataf(!\E_src1[26]~q ),
	.datag(gnd),
	.cin(\Add9~90 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~105_sumout ),
	.cout(\Add9~106 ),
	.shareout());
defparam \Add9~105 .extended_lut = "off";
defparam \Add9~105 .lut_mask = 64'h0000FF00000055AA;
defparam \Add9~105 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[26] (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\E_alu_result~17_combout ),
	.datac(!\Add9~105_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[26]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[26] .extended_lut = "off";
defparam \E_alu_result[26] .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \E_alu_result[26] .shared_arith = "off";

dffeas \M_alu_result[26] (
	.clk(clk_clk),
	.d(\E_alu_result[26]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_alu_result[26]~q ),
	.prn(vcc));
defparam \M_alu_result[26] .is_wysiwyg = "true";
defparam \M_alu_result[26] .power_up = "low";

cyclonev_lcell_comb \A_slow_inst_result_nxt[26]~24 (
	.dataa(!\A_ctrl_ld32~q ),
	.datab(!\A_ld_align_byte2_byte3_fill~q ),
	.datac(!src0_valid),
	.datad(!av_readdata_pre_26),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[26]~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[26]~24 .extended_lut = "off";
defparam \A_slow_inst_result_nxt[26]~24 .lut_mask = 64'h27FF27FF27FF27FF;
defparam \A_slow_inst_result_nxt[26]~24 .shared_arith = "off";

cyclonev_lcell_comb \A_slow_inst_result_nxt[26]~16 (
	.dataa(!\A_ctrl_ld32~q ),
	.datab(!\d_readdata_d1[26]~q ),
	.datac(!\A_slow_ld_data_fill_bit~0_combout ),
	.datad(!src0_valid1),
	.datae(!q_a_26),
	.dataf(!\A_slow_inst_result_nxt[26]~24_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[26]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[26]~16 .extended_lut = "off";
defparam \A_slow_inst_result_nxt[26]~16 .lut_mask = 64'h7FFFFFFFBFFFFFFF;
defparam \A_slow_inst_result_nxt[26]~16 .shared_arith = "off";

dffeas \A_slow_inst_result[26] (
	.clk(clk_clk),
	.d(\A_slow_inst_result_nxt[26]~16_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_ctrl_ld~q ),
	.q(\A_slow_inst_result[26]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[26] .is_wysiwyg = "true";
defparam \A_slow_inst_result[26] .power_up = "low";

cyclonev_lcell_comb \M_rot[2]~20 (
	.dataa(!\M_rot_prestep2[26]~q ),
	.datab(!\M_rot_prestep2[18]~q ),
	.datac(!\M_rot_prestep2[10]~q ),
	.datad(!\M_rot_prestep2[2]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[2]~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[2]~20 .extended_lut = "off";
defparam \M_rot[2]~20 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[2]~20 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~20 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_mask[2]~q ),
	.datac(!\M_rot_pass3~q ),
	.datad(!\M_rot_sel_fill3~q ),
	.datae(!\M_rot[2]~20_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~20 .extended_lut = "off";
defparam \A_shift_rot_result~20 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~20 .shared_arith = "off";

dffeas \A_shift_rot_result[26] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~20_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_shift_rot_result[26]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[26] .is_wysiwyg = "true";
defparam \A_shift_rot_result[26] .power_up = "low";

dffeas \A_inst_result[26] (
	.clk(clk_clk),
	.d(\M_alu_result[26]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\A_inst_result[26]~1_combout ),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_inst_result[26]~q ),
	.prn(vcc));
defparam \A_inst_result[26] .is_wysiwyg = "true";
defparam \A_inst_result[26] .power_up = "low";

cyclonev_lcell_comb \Add11~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[10]~q ),
	.datae(gnd),
	.dataf(!\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[26]~q ),
	.datag(gnd),
	.cin(\Add11~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add11~33_sumout ),
	.cout(\Add11~34 ),
	.shareout());
defparam \Add11~33 .extended_lut = "off";
defparam \Add11~33 .lut_mask = 64'h0000FF00000000FF;
defparam \Add11~33 .shared_arith = "off";

dffeas \A_mul_s1[10] (
	.clk(clk_clk),
	.d(\Add11~33_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_mul_s1[10]~q ),
	.prn(vcc));
defparam \A_mul_s1[10] .is_wysiwyg = "true";
defparam \A_mul_s1[10] .power_up = "low";

dffeas \A_mul_cell_p3[10] (
	.clk(clk_clk),
	.d(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p3|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[10]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_mul_cell_p3[10]~q ),
	.prn(vcc));
defparam \A_mul_cell_p3[10] .is_wysiwyg = "true";
defparam \A_mul_cell_p3[10] .power_up = "low";

cyclonev_lcell_comb \Add12~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_mul_s1[10]~q ),
	.datae(gnd),
	.dataf(!\A_mul_cell_p3[10]~q ),
	.datag(gnd),
	.cin(\Add12~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add12~33_sumout ),
	.cout(\Add12~34 ),
	.shareout());
defparam \Add12~33 .extended_lut = "off";
defparam \Add12~33 .lut_mask = 64'h0000FF00000000FF;
defparam \Add12~33 .shared_arith = "off";

cyclonev_lcell_comb \A_wr_data_unfiltered[26]~22 (
	.dataa(!\A_slow_inst_result[26]~q ),
	.datab(!\A_shift_rot_result[26]~q ),
	.datac(!\A_inst_result[26]~q ),
	.datad(!\Add12~33_sumout ),
	.datae(!\A_wr_data_unfiltered[15]~0_combout ),
	.dataf(!\A_wr_data_unfiltered[15]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[26]~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[26]~22 .extended_lut = "off";
defparam \A_wr_data_unfiltered[26]~22 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_wr_data_unfiltered[26]~22 .shared_arith = "off";

dffeas \W_wr_data[26] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[26]~22_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[26]~q ),
	.prn(vcc));
defparam \W_wr_data[26] .is_wysiwyg = "true";
defparam \W_wr_data[26] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[26]~19 (
	.dataa(!\M_alu_result[26]~q ),
	.datab(!\A_wr_data_unfiltered[26]~22_combout ),
	.datac(!\first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[26] ),
	.datad(!\W_wr_data[26]~q ),
	.datae(!\E_src1[26]~0_combout ),
	.dataf(!\E_src1[26]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[26]~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[26]~19 .extended_lut = "off";
defparam \D_src1_reg[26]~19 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[26]~19 .shared_arith = "off";

dffeas \E_src1[26] (
	.clk(clk_clk),
	.d(\D_src1_reg[26]~19_combout ),
	.asdata(\E_alu_result[26]~combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\Equal303~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(!\A_mem_stall~q ),
	.q(\E_src1[26]~q ),
	.prn(vcc));
defparam \E_src1[26] .is_wysiwyg = "true";
defparam \E_src1[26] .power_up = "low";

cyclonev_lcell_comb \E_alu_result~17 (
	.dataa(!\E_src2[26]~q ),
	.datab(!\E_src1[26]~q ),
	.datac(!\E_logic_op[1]~q ),
	.datad(!\E_logic_op[0]~q ),
	.datae(!\E_ctrl_logic~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result~17 .extended_lut = "off";
defparam \E_alu_result~17 .lut_mask = 64'h6996FFFF6996FFFF;
defparam \E_alu_result~17 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[26]~52 (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\D_src2_reg[0]~2_combout ),
	.datac(!\E_alu_result~17_combout ),
	.datad(!\Add9~105_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[26]~52_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[26]~52 .extended_lut = "off";
defparam \D_src2_reg[26]~52 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \D_src2_reg[26]~52 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[26]~53 (
	.dataa(!\D_src2_reg[0]~7_combout ),
	.datab(!\D_src2_reg[0]~8_combout ),
	.datac(!\D_src2_reg[0]~9_combout ),
	.datad(!\M_alu_result[26]~q ),
	.datae(!\A_wr_data_unfiltered[26]~22_combout ),
	.dataf(!\W_wr_data[26]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[26]~53_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[26]~53 .extended_lut = "off";
defparam \D_src2_reg[26]~53 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \D_src2_reg[26]~53 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[26]~17 (
	.dataa(!\D_iw[16]~q ),
	.datab(!\D_ctrl_hi_imm16~q ),
	.datac(!\D_iw[21]~q ),
	.datad(!\D_ctrl_unsigned_lo_imm16~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[26]~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[26]~17 .extended_lut = "off";
defparam \D_src2[26]~17 .lut_mask = 64'h7FDF7FDF7FDF7FDF;
defparam \D_src2[26]~17 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[26]~18 (
	.dataa(!\D_src2_reg[0]~6_combout ),
	.datab(!\D_ctrl_src2_choose_imm~q ),
	.datac(!\D_src2_reg[26]~52_combout ),
	.datad(!\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[26] ),
	.datae(!\D_src2_reg[26]~53_combout ),
	.dataf(!\D_src2[26]~17_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[26]~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[26]~18 .extended_lut = "off";
defparam \D_src2[26]~18 .lut_mask = 64'h47FFFFFFFFFFFFFF;
defparam \D_src2[26]~18 .shared_arith = "off";

dffeas \E_src2[26] (
	.clk(clk_clk),
	.d(\D_src2[26]~18_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src2[30]~1_combout ),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_src2[26]~q ),
	.prn(vcc));
defparam \E_src2[26] .is_wysiwyg = "true";
defparam \E_src2[26] .power_up = "low";

cyclonev_lcell_comb \Add9~101 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[27]~q ),
	.datae(gnd),
	.dataf(!\E_src1[27]~q ),
	.datag(gnd),
	.cin(\Add9~106 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~101_sumout ),
	.cout(\Add9~102 ),
	.shareout());
defparam \Add9~101 .extended_lut = "off";
defparam \Add9~101 .lut_mask = 64'h0000FF00000055AA;
defparam \Add9~101 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[27] (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\E_alu_result~14_combout ),
	.datac(!\Add9~101_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[27]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[27] .extended_lut = "off";
defparam \E_alu_result[27] .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \E_alu_result[27] .shared_arith = "off";

dffeas \M_alu_result[27] (
	.clk(clk_clk),
	.d(\E_alu_result[27]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_alu_result[27]~q ),
	.prn(vcc));
defparam \M_alu_result[27] .is_wysiwyg = "true";
defparam \M_alu_result[27] .power_up = "low";

cyclonev_lcell_comb \A_slow_inst_result_nxt[27]~25 (
	.dataa(!\A_ctrl_ld32~q ),
	.datab(!\A_ld_align_byte2_byte3_fill~q ),
	.datac(!src0_valid),
	.datad(!src_payload2),
	.datae(!av_readdata_pre_27),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[27]~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[27]~25 .extended_lut = "off";
defparam \A_slow_inst_result_nxt[27]~25 .lut_mask = 64'hFFFFFFD8FFFFFFD8;
defparam \A_slow_inst_result_nxt[27]~25 .shared_arith = "off";

cyclonev_lcell_comb \A_slow_inst_result_nxt[27]~15 (
	.dataa(!\A_ctrl_ld32~q ),
	.datab(!\d_readdata_d1[27]~q ),
	.datac(!\A_slow_ld_data_fill_bit~0_combout ),
	.datad(!src0_valid1),
	.datae(!q_a_27),
	.dataf(!\A_slow_inst_result_nxt[27]~25_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[27]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[27]~15 .extended_lut = "off";
defparam \A_slow_inst_result_nxt[27]~15 .lut_mask = 64'h7FFFFFFFBFFFFFFF;
defparam \A_slow_inst_result_nxt[27]~15 .shared_arith = "off";

dffeas \A_slow_inst_result[27] (
	.clk(clk_clk),
	.d(\A_slow_inst_result_nxt[27]~15_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_ctrl_ld~q ),
	.q(\A_slow_inst_result[27]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[27] .is_wysiwyg = "true";
defparam \A_slow_inst_result[27] .power_up = "low";

cyclonev_lcell_comb \M_rot[3]~17 (
	.dataa(!\M_rot_prestep2[27]~q ),
	.datab(!\M_rot_prestep2[19]~q ),
	.datac(!\M_rot_prestep2[11]~q ),
	.datad(!\M_rot_prestep2[3]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[3]~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[3]~17 .extended_lut = "off";
defparam \M_rot[3]~17 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[3]~17 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~17 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_mask[3]~q ),
	.datac(!\M_rot_pass3~q ),
	.datad(!\M_rot_sel_fill3~q ),
	.datae(!\M_rot[3]~17_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~17 .extended_lut = "off";
defparam \A_shift_rot_result~17 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~17 .shared_arith = "off";

dffeas \A_shift_rot_result[27] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~17_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_shift_rot_result[27]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[27] .is_wysiwyg = "true";
defparam \A_shift_rot_result[27] .power_up = "low";

dffeas \A_inst_result[27] (
	.clk(clk_clk),
	.d(\M_alu_result[27]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\A_inst_result[26]~1_combout ),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_inst_result[27]~q ),
	.prn(vcc));
defparam \A_inst_result[27] .is_wysiwyg = "true";
defparam \A_inst_result[27] .power_up = "low";

cyclonev_lcell_comb \Add11~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[11]~q ),
	.datae(gnd),
	.dataf(!\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[27]~q ),
	.datag(gnd),
	.cin(\Add11~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add11~29_sumout ),
	.cout(\Add11~30 ),
	.shareout());
defparam \Add11~29 .extended_lut = "off";
defparam \Add11~29 .lut_mask = 64'h0000FF00000000FF;
defparam \Add11~29 .shared_arith = "off";

dffeas \A_mul_s1[11] (
	.clk(clk_clk),
	.d(\Add11~29_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_mul_s1[11]~q ),
	.prn(vcc));
defparam \A_mul_s1[11] .is_wysiwyg = "true";
defparam \A_mul_s1[11] .power_up = "low";

dffeas \A_mul_cell_p3[11] (
	.clk(clk_clk),
	.d(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p3|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[11]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_mul_cell_p3[11]~q ),
	.prn(vcc));
defparam \A_mul_cell_p3[11] .is_wysiwyg = "true";
defparam \A_mul_cell_p3[11] .power_up = "low";

cyclonev_lcell_comb \Add12~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_mul_s1[11]~q ),
	.datae(gnd),
	.dataf(!\A_mul_cell_p3[11]~q ),
	.datag(gnd),
	.cin(\Add12~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add12~29_sumout ),
	.cout(\Add12~30 ),
	.shareout());
defparam \Add12~29 .extended_lut = "off";
defparam \Add12~29 .lut_mask = 64'h0000FF00000000FF;
defparam \Add12~29 .shared_arith = "off";

cyclonev_lcell_comb \A_wr_data_unfiltered[27]~19 (
	.dataa(!\A_slow_inst_result[27]~q ),
	.datab(!\A_shift_rot_result[27]~q ),
	.datac(!\A_inst_result[27]~q ),
	.datad(!\Add12~29_sumout ),
	.datae(!\A_wr_data_unfiltered[15]~0_combout ),
	.dataf(!\A_wr_data_unfiltered[15]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[27]~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[27]~19 .extended_lut = "off";
defparam \A_wr_data_unfiltered[27]~19 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_wr_data_unfiltered[27]~19 .shared_arith = "off";

dffeas \W_wr_data[27] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[27]~19_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[27]~q ),
	.prn(vcc));
defparam \W_wr_data[27] .is_wysiwyg = "true";
defparam \W_wr_data[27] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[27]~13 (
	.dataa(!\M_alu_result[27]~q ),
	.datab(!\A_wr_data_unfiltered[27]~19_combout ),
	.datac(!\first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[27] ),
	.datad(!\W_wr_data[27]~q ),
	.datae(!\E_src1[26]~0_combout ),
	.dataf(!\E_src1[26]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[27]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[27]~13 .extended_lut = "off";
defparam \D_src1_reg[27]~13 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[27]~13 .shared_arith = "off";

dffeas \E_src1[27] (
	.clk(clk_clk),
	.d(\D_src1_reg[27]~13_combout ),
	.asdata(\E_alu_result[27]~combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\Equal303~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(!\A_mem_stall~q ),
	.q(\E_src1[27]~q ),
	.prn(vcc));
defparam \E_src1[27] .is_wysiwyg = "true";
defparam \E_src1[27] .power_up = "low";

cyclonev_lcell_comb \E_alu_result~14 (
	.dataa(!\E_src2[27]~q ),
	.datab(!\E_src1[27]~q ),
	.datac(!\E_logic_op[1]~q ),
	.datad(!\E_logic_op[0]~q ),
	.datae(!\E_ctrl_logic~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result~14 .extended_lut = "off";
defparam \E_alu_result~14 .lut_mask = 64'h6996FFFF6996FFFF;
defparam \E_alu_result~14 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[27]~45 (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\D_src2_reg[0]~2_combout ),
	.datac(!\E_alu_result~14_combout ),
	.datad(!\Add9~101_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[27]~45_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[27]~45 .extended_lut = "off";
defparam \D_src2_reg[27]~45 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \D_src2_reg[27]~45 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[27]~34 (
	.dataa(!\D_src2_reg[0]~7_combout ),
	.datab(!\D_src2_reg[0]~8_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[27]~34_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[27]~34 .extended_lut = "off";
defparam \D_src2_reg[27]~34 .lut_mask = 64'h7777777777777777;
defparam \D_src2_reg[27]~34 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[27]~46 (
	.dataa(!\D_ctrl_b_is_dst~q ),
	.datab(!\A_regnum_b_cmp_D~q ),
	.datac(!\M_regnum_b_cmp_D~q ),
	.datad(!\M_alu_result[27]~q ),
	.datae(!\W_wr_data[27]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[27]~46_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[27]~46 .extended_lut = "off";
defparam \D_src2_reg[27]~46 .lut_mask = 64'hDEFFFFFFDEFFFFFF;
defparam \D_src2_reg[27]~46 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[27]~47 (
	.dataa(!\D_src2_reg[0]~9_combout ),
	.datab(!\A_wr_data_unfiltered[27]~19_combout ),
	.datac(!\D_src2_reg[27]~34_combout ),
	.datad(!\D_src2_reg[27]~46_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[27]~47_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[27]~47 .extended_lut = "off";
defparam \D_src2_reg[27]~47 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \D_src2_reg[27]~47 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[27]~14 (
	.dataa(!\D_ctrl_hi_imm16~q ),
	.datab(!\D_iw[21]~q ),
	.datac(!\D_ctrl_unsigned_lo_imm16~q ),
	.datad(!\D_iw[17]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[27]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[27]~14 .extended_lut = "off";
defparam \D_src2[27]~14 .lut_mask = 64'h7BFF7BFF7BFF7BFF;
defparam \D_src2[27]~14 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[27]~15 (
	.dataa(!\D_src2_reg[0]~6_combout ),
	.datab(!\D_ctrl_src2_choose_imm~q ),
	.datac(!\D_src2_reg[27]~45_combout ),
	.datad(!\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[27] ),
	.datae(!\D_src2_reg[27]~47_combout ),
	.dataf(!\D_src2[27]~14_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[27]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[27]~15 .extended_lut = "off";
defparam \D_src2[27]~15 .lut_mask = 64'h47FFFFFFFFFFFFFF;
defparam \D_src2[27]~15 .shared_arith = "off";

dffeas \E_src2[27] (
	.clk(clk_clk),
	.d(\D_src2[27]~15_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src2[30]~1_combout ),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_src2[27]~q ),
	.prn(vcc));
defparam \E_src2[27] .is_wysiwyg = "true";
defparam \E_src2[27] .power_up = "low";

cyclonev_lcell_comb \Add9~97 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[28]~q ),
	.datae(gnd),
	.dataf(!\E_src1[28]~q ),
	.datag(gnd),
	.cin(\Add9~102 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~97_sumout ),
	.cout(\Add9~98 ),
	.shareout());
defparam \Add9~97 .extended_lut = "off";
defparam \Add9~97 .lut_mask = 64'h0000FF00000055AA;
defparam \Add9~97 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[28] (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\E_alu_result~12_combout ),
	.datac(!\Add9~97_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[28]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[28] .extended_lut = "off";
defparam \E_alu_result[28] .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \E_alu_result[28] .shared_arith = "off";

dffeas \M_alu_result[28] (
	.clk(clk_clk),
	.d(\E_alu_result[28]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_alu_result[28]~q ),
	.prn(vcc));
defparam \M_alu_result[28] .is_wysiwyg = "true";
defparam \M_alu_result[28] .power_up = "low";

cyclonev_lcell_comb \A_slow_inst_result_nxt[28]~26 (
	.dataa(!\A_ctrl_ld32~q ),
	.datab(!\A_ld_align_byte2_byte3_fill~q ),
	.datac(!src0_valid),
	.datad(!src_payload2),
	.datae(!av_readdata_pre_28),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[28]~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[28]~26 .extended_lut = "off";
defparam \A_slow_inst_result_nxt[28]~26 .lut_mask = 64'hFFFFFFD8FFFFFFD8;
defparam \A_slow_inst_result_nxt[28]~26 .shared_arith = "off";

cyclonev_lcell_comb \A_slow_inst_result_nxt[28]~14 (
	.dataa(!\A_ctrl_ld32~q ),
	.datab(!\d_readdata_d1[28]~q ),
	.datac(!\A_slow_ld_data_fill_bit~0_combout ),
	.datad(!src0_valid1),
	.datae(!q_a_28),
	.dataf(!\A_slow_inst_result_nxt[28]~26_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[28]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[28]~14 .extended_lut = "off";
defparam \A_slow_inst_result_nxt[28]~14 .lut_mask = 64'h7FFFFFFFBFFFFFFF;
defparam \A_slow_inst_result_nxt[28]~14 .shared_arith = "off";

dffeas \A_slow_inst_result[28] (
	.clk(clk_clk),
	.d(\A_slow_inst_result_nxt[28]~14_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_ctrl_ld~q ),
	.q(\A_slow_inst_result[28]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[28] .is_wysiwyg = "true";
defparam \A_slow_inst_result[28] .power_up = "low";

cyclonev_lcell_comb \M_rot[4]~15 (
	.dataa(!\M_rot_prestep2[28]~q ),
	.datab(!\M_rot_prestep2[20]~q ),
	.datac(!\M_rot_prestep2[12]~q ),
	.datad(!\M_rot_prestep2[4]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[4]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[4]~15 .extended_lut = "off";
defparam \M_rot[4]~15 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[4]~15 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~15 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_mask[4]~q ),
	.datac(!\M_rot_pass3~q ),
	.datad(!\M_rot_sel_fill3~q ),
	.datae(!\M_rot[4]~15_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~15 .extended_lut = "off";
defparam \A_shift_rot_result~15 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~15 .shared_arith = "off";

dffeas \A_shift_rot_result[28] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~15_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_shift_rot_result[28]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[28] .is_wysiwyg = "true";
defparam \A_shift_rot_result[28] .power_up = "low";

dffeas \A_inst_result[28] (
	.clk(clk_clk),
	.d(\M_alu_result[28]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\A_inst_result[26]~1_combout ),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_inst_result[28]~q ),
	.prn(vcc));
defparam \A_inst_result[28] .is_wysiwyg = "true";
defparam \A_inst_result[28] .power_up = "low";

cyclonev_lcell_comb \Add11~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[12]~q ),
	.datae(gnd),
	.dataf(!\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[28]~q ),
	.datag(gnd),
	.cin(\Add11~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add11~25_sumout ),
	.cout(\Add11~26 ),
	.shareout());
defparam \Add11~25 .extended_lut = "off";
defparam \Add11~25 .lut_mask = 64'h0000FF00000000FF;
defparam \Add11~25 .shared_arith = "off";

dffeas \A_mul_s1[12] (
	.clk(clk_clk),
	.d(\Add11~25_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_mul_s1[12]~q ),
	.prn(vcc));
defparam \A_mul_s1[12] .is_wysiwyg = "true";
defparam \A_mul_s1[12] .power_up = "low";

dffeas \A_mul_cell_p3[12] (
	.clk(clk_clk),
	.d(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p3|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[12]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_mul_cell_p3[12]~q ),
	.prn(vcc));
defparam \A_mul_cell_p3[12] .is_wysiwyg = "true";
defparam \A_mul_cell_p3[12] .power_up = "low";

cyclonev_lcell_comb \Add12~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_mul_s1[12]~q ),
	.datae(gnd),
	.dataf(!\A_mul_cell_p3[12]~q ),
	.datag(gnd),
	.cin(\Add12~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add12~25_sumout ),
	.cout(\Add12~26 ),
	.shareout());
defparam \Add12~25 .extended_lut = "off";
defparam \Add12~25 .lut_mask = 64'h0000FF00000000FF;
defparam \Add12~25 .shared_arith = "off";

cyclonev_lcell_comb \A_wr_data_unfiltered[28]~17 (
	.dataa(!\A_slow_inst_result[28]~q ),
	.datab(!\A_shift_rot_result[28]~q ),
	.datac(!\A_inst_result[28]~q ),
	.datad(!\Add12~25_sumout ),
	.datae(!\A_wr_data_unfiltered[15]~0_combout ),
	.dataf(!\A_wr_data_unfiltered[15]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[28]~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[28]~17 .extended_lut = "off";
defparam \A_wr_data_unfiltered[28]~17 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_wr_data_unfiltered[28]~17 .shared_arith = "off";

dffeas \W_wr_data[28] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[28]~17_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[28]~q ),
	.prn(vcc));
defparam \W_wr_data[28] .is_wysiwyg = "true";
defparam \W_wr_data[28] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[28]~11 (
	.dataa(!\M_alu_result[28]~q ),
	.datab(!\A_wr_data_unfiltered[28]~17_combout ),
	.datac(!\first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[28] ),
	.datad(!\W_wr_data[28]~q ),
	.datae(!\E_src1[26]~0_combout ),
	.dataf(!\E_src1[26]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[28]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[28]~11 .extended_lut = "off";
defparam \D_src1_reg[28]~11 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[28]~11 .shared_arith = "off";

dffeas \E_src1[28] (
	.clk(clk_clk),
	.d(\D_src1_reg[28]~11_combout ),
	.asdata(\E_alu_result[28]~combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\Equal303~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(!\A_mem_stall~q ),
	.q(\E_src1[28]~q ),
	.prn(vcc));
defparam \E_src1[28] .is_wysiwyg = "true";
defparam \E_src1[28] .power_up = "low";

cyclonev_lcell_comb \E_alu_result~12 (
	.dataa(!\E_src2[28]~q ),
	.datab(!\E_src1[28]~q ),
	.datac(!\E_logic_op[1]~q ),
	.datad(!\E_logic_op[0]~q ),
	.datae(!\E_ctrl_logic~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result~12 .extended_lut = "off";
defparam \E_alu_result~12 .lut_mask = 64'h6996FFFF6996FFFF;
defparam \E_alu_result~12 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[28]~40 (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\D_src2_reg[0]~2_combout ),
	.datac(!\E_alu_result~12_combout ),
	.datad(!\Add9~97_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[28]~40_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[28]~40 .extended_lut = "off";
defparam \D_src2_reg[28]~40 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \D_src2_reg[28]~40 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[28]~41 (
	.dataa(!\D_ctrl_b_is_dst~q ),
	.datab(!\A_regnum_b_cmp_D~q ),
	.datac(!\M_regnum_b_cmp_D~q ),
	.datad(!\M_alu_result[28]~q ),
	.datae(!\W_wr_data[28]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[28]~41_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[28]~41 .extended_lut = "off";
defparam \D_src2_reg[28]~41 .lut_mask = 64'hDEFFFFFFDEFFFFFF;
defparam \D_src2_reg[28]~41 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[28]~42 (
	.dataa(!\D_src2_reg[0]~9_combout ),
	.datab(!\D_src2_reg[27]~34_combout ),
	.datac(!\A_wr_data_unfiltered[28]~17_combout ),
	.datad(!\D_src2_reg[28]~41_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[28]~42_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[28]~42 .extended_lut = "off";
defparam \D_src2_reg[28]~42 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \D_src2_reg[28]~42 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[28]~12 (
	.dataa(!\D_ctrl_hi_imm16~q ),
	.datab(!\D_iw[21]~q ),
	.datac(!\D_ctrl_unsigned_lo_imm16~q ),
	.datad(!\D_iw[18]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[28]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[28]~12 .extended_lut = "off";
defparam \D_src2[28]~12 .lut_mask = 64'h7BFF7BFF7BFF7BFF;
defparam \D_src2[28]~12 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[28]~13 (
	.dataa(!\D_src2_reg[0]~6_combout ),
	.datab(!\D_ctrl_src2_choose_imm~q ),
	.datac(!\D_src2_reg[28]~40_combout ),
	.datad(!\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[28] ),
	.datae(!\D_src2_reg[28]~42_combout ),
	.dataf(!\D_src2[28]~12_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[28]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[28]~13 .extended_lut = "off";
defparam \D_src2[28]~13 .lut_mask = 64'h47FFFFFFFFFFFFFF;
defparam \D_src2[28]~13 .shared_arith = "off";

dffeas \E_src2[28] (
	.clk(clk_clk),
	.d(\D_src2[28]~13_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src2[30]~1_combout ),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_src2[28]~q ),
	.prn(vcc));
defparam \E_src2[28] .is_wysiwyg = "true";
defparam \E_src2[28] .power_up = "low";

cyclonev_lcell_comb \Add9~129 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[29]~q ),
	.datae(gnd),
	.dataf(!\E_src1[29]~q ),
	.datag(gnd),
	.cin(\Add9~98 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~129_sumout ),
	.cout(\Add9~130 ),
	.shareout());
defparam \Add9~129 .extended_lut = "off";
defparam \Add9~129 .lut_mask = 64'h0000FF00000055AA;
defparam \Add9~129 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[29] (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\E_alu_result~24_combout ),
	.datac(!\Add9~129_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[29]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[29] .extended_lut = "off";
defparam \E_alu_result[29] .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \E_alu_result[29] .shared_arith = "off";

dffeas \M_alu_result[29] (
	.clk(clk_clk),
	.d(\E_alu_result[29]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_alu_result[29]~q ),
	.prn(vcc));
defparam \M_alu_result[29] .is_wysiwyg = "true";
defparam \M_alu_result[29] .power_up = "low";

cyclonev_lcell_comb \A_slow_inst_result_nxt[29]~28 (
	.dataa(!\A_ctrl_ld32~q ),
	.datab(!\A_ld_align_byte2_byte3_fill~q ),
	.datac(!src0_valid),
	.datad(!av_readdata_pre_29),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[29]~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[29]~28 .extended_lut = "off";
defparam \A_slow_inst_result_nxt[29]~28 .lut_mask = 64'h27FF27FF27FF27FF;
defparam \A_slow_inst_result_nxt[29]~28 .shared_arith = "off";

cyclonev_lcell_comb \A_slow_inst_result_nxt[29]~23 (
	.dataa(!\A_ctrl_ld32~q ),
	.datab(!\d_readdata_d1[29]~q ),
	.datac(!\A_slow_ld_data_fill_bit~0_combout ),
	.datad(!src0_valid1),
	.datae(!q_a_29),
	.dataf(!\A_slow_inst_result_nxt[29]~28_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[29]~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[29]~23 .extended_lut = "off";
defparam \A_slow_inst_result_nxt[29]~23 .lut_mask = 64'h7FFFFFFFBFFFFFFF;
defparam \A_slow_inst_result_nxt[29]~23 .shared_arith = "off";

dffeas \A_slow_inst_result[29] (
	.clk(clk_clk),
	.d(\A_slow_inst_result_nxt[29]~23_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_ctrl_ld~q ),
	.q(\A_slow_inst_result[29]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[29] .is_wysiwyg = "true";
defparam \A_slow_inst_result[29] .power_up = "low";

cyclonev_lcell_comb \M_rot[5]~31 (
	.dataa(!\M_rot_prestep2[29]~q ),
	.datab(!\M_rot_prestep2[21]~q ),
	.datac(!\M_rot_prestep2[13]~q ),
	.datad(!\M_rot_prestep2[5]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[5]~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[5]~31 .extended_lut = "off";
defparam \M_rot[5]~31 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[5]~31 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~31 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_mask[5]~q ),
	.datac(!\M_rot_pass3~q ),
	.datad(!\M_rot_sel_fill3~q ),
	.datae(!\M_rot[5]~31_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~31 .extended_lut = "off";
defparam \A_shift_rot_result~31 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~31 .shared_arith = "off";

dffeas \A_shift_rot_result[29] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~31_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_shift_rot_result[29]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[29] .is_wysiwyg = "true";
defparam \A_shift_rot_result[29] .power_up = "low";

dffeas \A_inst_result[29] (
	.clk(clk_clk),
	.d(\M_alu_result[29]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\A_inst_result[26]~1_combout ),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_inst_result[29]~q ),
	.prn(vcc));
defparam \A_inst_result[29] .is_wysiwyg = "true";
defparam \A_inst_result[29] .power_up = "low";

cyclonev_lcell_comb \Add11~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[13]~q ),
	.datae(gnd),
	.dataf(!\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[29]~q ),
	.datag(gnd),
	.cin(\Add11~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add11~61_sumout ),
	.cout(\Add11~62 ),
	.shareout());
defparam \Add11~61 .extended_lut = "off";
defparam \Add11~61 .lut_mask = 64'h0000FF00000000FF;
defparam \Add11~61 .shared_arith = "off";

dffeas \A_mul_s1[13] (
	.clk(clk_clk),
	.d(\Add11~61_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_mul_s1[13]~q ),
	.prn(vcc));
defparam \A_mul_s1[13] .is_wysiwyg = "true";
defparam \A_mul_s1[13] .power_up = "low";

dffeas \A_mul_cell_p3[13] (
	.clk(clk_clk),
	.d(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p3|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[13]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_mul_cell_p3[13]~q ),
	.prn(vcc));
defparam \A_mul_cell_p3[13] .is_wysiwyg = "true";
defparam \A_mul_cell_p3[13] .power_up = "low";

cyclonev_lcell_comb \Add12~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_mul_s1[13]~q ),
	.datae(gnd),
	.dataf(!\A_mul_cell_p3[13]~q ),
	.datag(gnd),
	.cin(\Add12~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add12~61_sumout ),
	.cout(\Add12~62 ),
	.shareout());
defparam \Add12~61 .extended_lut = "off";
defparam \Add12~61 .lut_mask = 64'h0000FF00000000FF;
defparam \Add12~61 .shared_arith = "off";

cyclonev_lcell_comb \A_wr_data_unfiltered[29]~33 (
	.dataa(!\A_slow_inst_result[29]~q ),
	.datab(!\A_shift_rot_result[29]~q ),
	.datac(!\A_inst_result[29]~q ),
	.datad(!\Add12~61_sumout ),
	.datae(!\A_wr_data_unfiltered[15]~0_combout ),
	.dataf(!\A_wr_data_unfiltered[15]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[29]~33_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[29]~33 .extended_lut = "off";
defparam \A_wr_data_unfiltered[29]~33 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_wr_data_unfiltered[29]~33 .shared_arith = "off";

dffeas \W_wr_data[29] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[29]~33_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[29]~q ),
	.prn(vcc));
defparam \W_wr_data[29] .is_wysiwyg = "true";
defparam \W_wr_data[29] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[29]~31 (
	.dataa(!\M_alu_result[29]~q ),
	.datab(!\A_wr_data_unfiltered[29]~33_combout ),
	.datac(!\first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[29] ),
	.datad(!\W_wr_data[29]~q ),
	.datae(!\E_src1[26]~0_combout ),
	.dataf(!\E_src1[26]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[29]~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[29]~31 .extended_lut = "off";
defparam \D_src1_reg[29]~31 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[29]~31 .shared_arith = "off";

dffeas \E_src1[29] (
	.clk(clk_clk),
	.d(\D_src1_reg[29]~31_combout ),
	.asdata(\E_alu_result[29]~combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\Equal303~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(!\A_mem_stall~q ),
	.q(\E_src1[29]~q ),
	.prn(vcc));
defparam \E_src1[29] .is_wysiwyg = "true";
defparam \E_src1[29] .power_up = "low";

cyclonev_lcell_comb \E_alu_result~24 (
	.dataa(!\E_src2[29]~q ),
	.datab(!\E_src1[29]~q ),
	.datac(!\E_logic_op[1]~q ),
	.datad(!\E_logic_op[0]~q ),
	.datae(!\E_ctrl_logic~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result~24 .extended_lut = "off";
defparam \E_alu_result~24 .lut_mask = 64'h6996FFFF6996FFFF;
defparam \E_alu_result~24 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[29]~70 (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\D_src2_reg[0]~2_combout ),
	.datac(!\E_alu_result~24_combout ),
	.datad(!\Add9~129_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[29]~70_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[29]~70 .extended_lut = "off";
defparam \D_src2_reg[29]~70 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \D_src2_reg[29]~70 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[29]~71 (
	.dataa(!\D_ctrl_b_is_dst~q ),
	.datab(!\A_regnum_b_cmp_D~q ),
	.datac(!\M_regnum_b_cmp_D~q ),
	.datad(!\M_alu_result[29]~q ),
	.datae(!\W_wr_data[29]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[29]~71_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[29]~71 .extended_lut = "off";
defparam \D_src2_reg[29]~71 .lut_mask = 64'hDEFFFFFFDEFFFFFF;
defparam \D_src2_reg[29]~71 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[29]~72 (
	.dataa(!\D_src2_reg[0]~9_combout ),
	.datab(!\D_src2_reg[27]~34_combout ),
	.datac(!\A_wr_data_unfiltered[29]~33_combout ),
	.datad(!\D_src2_reg[29]~71_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[29]~72_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[29]~72 .extended_lut = "off";
defparam \D_src2_reg[29]~72 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \D_src2_reg[29]~72 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[29]~27 (
	.dataa(!\D_ctrl_hi_imm16~q ),
	.datab(!\D_iw[21]~q ),
	.datac(!\D_ctrl_unsigned_lo_imm16~q ),
	.datad(!\D_iw[19]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[29]~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[29]~27 .extended_lut = "off";
defparam \D_src2[29]~27 .lut_mask = 64'h7BFF7BFF7BFF7BFF;
defparam \D_src2[29]~27 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[29]~28 (
	.dataa(!\D_src2_reg[0]~6_combout ),
	.datab(!\D_ctrl_src2_choose_imm~q ),
	.datac(!\D_src2_reg[29]~70_combout ),
	.datad(!\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[29] ),
	.datae(!\D_src2_reg[29]~72_combout ),
	.dataf(!\D_src2[29]~27_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[29]~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[29]~28 .extended_lut = "off";
defparam \D_src2[29]~28 .lut_mask = 64'h47FFFFFFFFFFFFFF;
defparam \D_src2[29]~28 .shared_arith = "off";

dffeas \E_src2[29] (
	.clk(clk_clk),
	.d(\D_src2[29]~28_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src2[30]~1_combout ),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_src2[29]~q ),
	.prn(vcc));
defparam \E_src2[29] .is_wysiwyg = "true";
defparam \E_src2[29] .power_up = "low";

cyclonev_lcell_comb \Add9~121 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[30]~q ),
	.datae(gnd),
	.dataf(!\E_src1[30]~q ),
	.datag(gnd),
	.cin(\Add9~130 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~121_sumout ),
	.cout(\Add9~122 ),
	.shareout());
defparam \Add9~121 .extended_lut = "off";
defparam \Add9~121 .lut_mask = 64'h0000FF00000055AA;
defparam \Add9~121 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[30]~57 (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\D_src2_reg[0]~2_combout ),
	.datac(!\E_alu_result~18_combout ),
	.datad(!\Add9~121_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[30]~57_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[30]~57 .extended_lut = "off";
defparam \D_src2_reg[30]~57 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \D_src2_reg[30]~57 .shared_arith = "off";

cyclonev_lcell_comb \A_slow_inst_result_nxt[30]~31 (
	.dataa(!\A_ctrl_ld32~q ),
	.datab(!\A_ld_align_byte2_byte3_fill~q ),
	.datac(!src0_valid),
	.datad(!src_payload2),
	.datae(!av_readdata_pre_30),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[30]~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[30]~31 .extended_lut = "off";
defparam \A_slow_inst_result_nxt[30]~31 .lut_mask = 64'hFFFFFFD8FFFFFFD8;
defparam \A_slow_inst_result_nxt[30]~31 .shared_arith = "off";

cyclonev_lcell_comb \A_slow_inst_result_nxt[30]~20 (
	.dataa(!\A_ctrl_ld32~q ),
	.datab(!\d_readdata_d1[30]~q ),
	.datac(!\A_slow_ld_data_fill_bit~0_combout ),
	.datad(!src0_valid1),
	.datae(!q_a_30),
	.dataf(!\A_slow_inst_result_nxt[30]~31_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[30]~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[30]~20 .extended_lut = "off";
defparam \A_slow_inst_result_nxt[30]~20 .lut_mask = 64'h7FFFFFFFBFFFFFFF;
defparam \A_slow_inst_result_nxt[30]~20 .shared_arith = "off";

dffeas \A_slow_inst_result[30] (
	.clk(clk_clk),
	.d(\A_slow_inst_result_nxt[30]~20_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_ctrl_ld~q ),
	.q(\A_slow_inst_result[30]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[30] .is_wysiwyg = "true";
defparam \A_slow_inst_result[30] .power_up = "low";

cyclonev_lcell_comb \M_rot[6]~24 (
	.dataa(!\M_rot_prestep2[30]~q ),
	.datab(!\M_rot_prestep2[22]~q ),
	.datac(!\M_rot_prestep2[14]~q ),
	.datad(!\M_rot_prestep2[6]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[6]~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[6]~24 .extended_lut = "off";
defparam \M_rot[6]~24 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[6]~24 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~24 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_mask[6]~q ),
	.datac(!\M_rot_pass3~q ),
	.datad(!\M_rot_sel_fill3~q ),
	.datae(!\M_rot[6]~24_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~24 .extended_lut = "off";
defparam \A_shift_rot_result~24 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~24 .shared_arith = "off";

dffeas \A_shift_rot_result[30] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~24_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_shift_rot_result[30]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[30] .is_wysiwyg = "true";
defparam \A_shift_rot_result[30] .power_up = "low";

dffeas \A_inst_result[30] (
	.clk(clk_clk),
	.d(\M_alu_result[30]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\A_inst_result[26]~1_combout ),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_inst_result[30]~q ),
	.prn(vcc));
defparam \A_inst_result[30] .is_wysiwyg = "true";
defparam \A_inst_result[30] .power_up = "low";

cyclonev_lcell_comb \Add11~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[14]~q ),
	.datae(gnd),
	.dataf(!\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[30]~q ),
	.datag(gnd),
	.cin(\Add11~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add11~49_sumout ),
	.cout(\Add11~50 ),
	.shareout());
defparam \Add11~49 .extended_lut = "off";
defparam \Add11~49 .lut_mask = 64'h0000FF00000000FF;
defparam \Add11~49 .shared_arith = "off";

dffeas \A_mul_s1[14] (
	.clk(clk_clk),
	.d(\Add11~49_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_mul_s1[14]~q ),
	.prn(vcc));
defparam \A_mul_s1[14] .is_wysiwyg = "true";
defparam \A_mul_s1[14] .power_up = "low";

dffeas \A_mul_cell_p3[14] (
	.clk(clk_clk),
	.d(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p3|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[14]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_mul_cell_p3[14]~q ),
	.prn(vcc));
defparam \A_mul_cell_p3[14] .is_wysiwyg = "true";
defparam \A_mul_cell_p3[14] .power_up = "low";

cyclonev_lcell_comb \Add12~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_mul_s1[14]~q ),
	.datae(gnd),
	.dataf(!\A_mul_cell_p3[14]~q ),
	.datag(gnd),
	.cin(\Add12~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add12~49_sumout ),
	.cout(\Add12~50 ),
	.shareout());
defparam \Add12~49 .extended_lut = "off";
defparam \Add12~49 .lut_mask = 64'h0000FF00000000FF;
defparam \Add12~49 .shared_arith = "off";

cyclonev_lcell_comb \A_wr_data_unfiltered[30]~26 (
	.dataa(!\A_slow_inst_result[30]~q ),
	.datab(!\A_shift_rot_result[30]~q ),
	.datac(!\A_inst_result[30]~q ),
	.datad(!\Add12~49_sumout ),
	.datae(!\A_wr_data_unfiltered[15]~0_combout ),
	.dataf(!\A_wr_data_unfiltered[15]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[30]~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[30]~26 .extended_lut = "off";
defparam \A_wr_data_unfiltered[30]~26 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_wr_data_unfiltered[30]~26 .shared_arith = "off";

dffeas \W_wr_data[30] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[30]~26_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[30]~q ),
	.prn(vcc));
defparam \W_wr_data[30] .is_wysiwyg = "true";
defparam \W_wr_data[30] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[30]~58 (
	.dataa(!\D_ctrl_b_is_dst~q ),
	.datab(!\A_regnum_b_cmp_D~q ),
	.datac(!\M_regnum_b_cmp_D~q ),
	.datad(!\M_alu_result[30]~q ),
	.datae(!\W_wr_data[30]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[30]~58_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[30]~58 .extended_lut = "off";
defparam \D_src2_reg[30]~58 .lut_mask = 64'hDEFFFFFFDEFFFFFF;
defparam \D_src2_reg[30]~58 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[30]~59 (
	.dataa(!\D_src2_reg[0]~9_combout ),
	.datab(!\D_src2_reg[27]~34_combout ),
	.datac(!\A_wr_data_unfiltered[30]~26_combout ),
	.datad(!\D_src2_reg[30]~58_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[30]~59_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[30]~59 .extended_lut = "off";
defparam \D_src2_reg[30]~59 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \D_src2_reg[30]~59 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[30]~22 (
	.dataa(!\D_ctrl_hi_imm16~q ),
	.datab(!\D_iw[21]~q ),
	.datac(!\D_ctrl_unsigned_lo_imm16~q ),
	.datad(!\D_iw[20]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[30]~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[30]~22 .extended_lut = "off";
defparam \D_src2[30]~22 .lut_mask = 64'h7BFF7BFF7BFF7BFF;
defparam \D_src2[30]~22 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[30]~23 (
	.dataa(!\D_src2_reg[0]~6_combout ),
	.datab(!\D_ctrl_src2_choose_imm~q ),
	.datac(!\D_src2_reg[30]~57_combout ),
	.datad(!\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[30] ),
	.datae(!\D_src2_reg[30]~59_combout ),
	.dataf(!\D_src2[30]~22_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[30]~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[30]~23 .extended_lut = "off";
defparam \D_src2[30]~23 .lut_mask = 64'h47FFFFFFFFFFFFFF;
defparam \D_src2[30]~23 .shared_arith = "off";

dffeas \E_src2[30] (
	.clk(clk_clk),
	.d(\D_src2[30]~23_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src2[30]~1_combout ),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_src2[30]~q ),
	.prn(vcc));
defparam \E_src2[30] .is_wysiwyg = "true";
defparam \E_src2[30] .power_up = "low";

cyclonev_lcell_comb \E_logic_result[30]~5 (
	.dataa(!\E_src2[30]~q ),
	.datab(!\E_src1[30]~q ),
	.datac(!\E_logic_op[1]~q ),
	.datad(!\E_logic_op[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[30]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[30]~5 .extended_lut = "off";
defparam \E_logic_result[30]~5 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[30]~5 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result~18 (
	.dataa(!\E_logic_result[30]~5_combout ),
	.datab(!\E_ctrl_logic~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result~18 .extended_lut = "off";
defparam \E_alu_result~18 .lut_mask = 64'h7777777777777777;
defparam \E_alu_result~18 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[30] (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\E_alu_result~18_combout ),
	.datac(!\Add9~121_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[30]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[30] .extended_lut = "off";
defparam \E_alu_result[30] .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \E_alu_result[30] .shared_arith = "off";

dffeas \M_alu_result[30] (
	.clk(clk_clk),
	.d(\E_alu_result[30]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_alu_result[30]~q ),
	.prn(vcc));
defparam \M_alu_result[30] .is_wysiwyg = "true";
defparam \M_alu_result[30] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[30]~23 (
	.dataa(!\M_alu_result[30]~q ),
	.datab(!\A_wr_data_unfiltered[30]~26_combout ),
	.datac(!\first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[30] ),
	.datad(!\W_wr_data[30]~q ),
	.datae(!\E_src1[26]~0_combout ),
	.dataf(!\E_src1[26]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[30]~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[30]~23 .extended_lut = "off";
defparam \D_src1_reg[30]~23 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[30]~23 .shared_arith = "off";

dffeas \E_src1[30] (
	.clk(clk_clk),
	.d(\D_src1_reg[30]~23_combout ),
	.asdata(\E_alu_result[30]~combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\Equal303~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(!\A_mem_stall~q ),
	.q(\E_src1[30]~q ),
	.prn(vcc));
defparam \E_src1[30] .is_wysiwyg = "true";
defparam \E_src1[30] .power_up = "low";

cyclonev_lcell_comb \E_rot_step1[30]~16 (
	.dataa(!\E_src1[30]~q ),
	.datab(!\E_src1[29]~q ),
	.datac(!\E_src1[28]~q ),
	.datad(!\E_src1[27]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add10~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[30]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[30]~16 .extended_lut = "off";
defparam \E_rot_step1[30]~16 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[30]~16 .shared_arith = "off";

dffeas \M_rot_prestep2[2] (
	.clk(clk_clk),
	.d(\E_rot_step1[30]~16_combout ),
	.asdata(\E_rot_step1[2]~17_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add10~1_combout ),
	.ena(!\A_mem_stall~q ),
	.q(\M_rot_prestep2[2]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[2] .is_wysiwyg = "true";
defparam \M_rot_prestep2[2] .power_up = "low";

cyclonev_lcell_comb \M_rot[2]~2 (
	.dataa(!\M_rot_prestep2[2]~q ),
	.datab(!\M_rot_prestep2[26]~q ),
	.datac(!\M_rot_prestep2[18]~q ),
	.datad(!\M_rot_prestep2[10]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[2]~2 .extended_lut = "off";
defparam \M_rot[2]~2 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[2]~2 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~2 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_pass0~q ),
	.datac(!\M_rot_sel_fill0~q ),
	.datad(!\M_rot_mask[2]~q ),
	.datae(!\M_rot[2]~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~2 .extended_lut = "off";
defparam \A_shift_rot_result~2 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~2 .shared_arith = "off";

dffeas \A_shift_rot_result[2] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_shift_rot_result[2]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[2] .is_wysiwyg = "true";
defparam \A_shift_rot_result[2] .power_up = "low";

cyclonev_lcell_comb \Equal327~0 (
	.dataa(!\E_iw[9]~q ),
	.datab(!\E_iw[7]~q ),
	.datac(!\E_iw[6]~q ),
	.datad(!\E_iw[10]~q ),
	.datae(!\E_iw[8]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal327~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal327~0 .extended_lut = "off";
defparam \Equal327~0 .lut_mask = 64'hFFBFFFFFFFBFFFFF;
defparam \Equal327~0 .shared_arith = "off";

cyclonev_lcell_comb \latched_oci_tb_hbreak_req_next~0 (
	.dataa(!W_debug_mode1),
	.datab(!\latched_oci_tb_hbreak_req~q ),
	.datac(!\hbreak_req~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\latched_oci_tb_hbreak_req_next~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \latched_oci_tb_hbreak_req_next~0 .extended_lut = "off";
defparam \latched_oci_tb_hbreak_req_next~0 .lut_mask = 64'h8B8B8B8B8B8B8B8B;
defparam \latched_oci_tb_hbreak_req_next~0 .shared_arith = "off";

dffeas latched_oci_tb_hbreak_req(
	.clk(clk_clk),
	.d(\latched_oci_tb_hbreak_req_next~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\latched_oci_tb_hbreak_req~q ),
	.prn(vcc));
defparam latched_oci_tb_hbreak_req.is_wysiwyg = "true";
defparam latched_oci_tb_hbreak_req.power_up = "low";

cyclonev_lcell_comb \A_exc_norm_intr_pri5_nxt~0 (
	.dataa(!\M_norm_intr_req~q ),
	.datab(!W_debug_mode1),
	.datac(!\the_first_nios2_system_cpu_cpu_nios2_oci|the_first_nios2_system_cpu_cpu_nios2_avalon_reg|oci_single_step_mode~q ),
	.datad(!\wait_for_one_post_bret_inst~0_combout ),
	.datae(!\latched_oci_tb_hbreak_req~q ),
	.dataf(!\the_first_nios2_system_cpu_cpu_nios2_oci|the_first_nios2_system_cpu_cpu_nios2_oci_debug|jtag_break~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_exc_norm_intr_pri5_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_exc_norm_intr_pri5_nxt~0 .extended_lut = "off";
defparam \A_exc_norm_intr_pri5_nxt~0 .lut_mask = 64'hFFFFFFFFFFFF7FFF;
defparam \A_exc_norm_intr_pri5_nxt~0 .shared_arith = "off";

dffeas A_exc_norm_intr_pri5(
	.clk(clk_clk),
	.d(\A_exc_norm_intr_pri5_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_exc_norm_intr_pri5~q ),
	.prn(vcc));
defparam A_exc_norm_intr_pri5.is_wysiwyg = "true";
defparam A_exc_norm_intr_pri5.power_up = "low";

cyclonev_lcell_comb \A_exc_trap_inst_pri15_nxt~0 (
	.dataa(!\M_exc_trap_inst_pri15~q ),
	.datab(!\M_norm_intr_req~q ),
	.datac(!\hbreak_req~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_exc_trap_inst_pri15_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_exc_trap_inst_pri15_nxt~0 .extended_lut = "off";
defparam \A_exc_trap_inst_pri15_nxt~0 .lut_mask = 64'hFDFDFDFDFDFDFDFD;
defparam \A_exc_trap_inst_pri15_nxt~0 .shared_arith = "off";

dffeas A_exc_trap_inst_pri15(
	.clk(clk_clk),
	.d(\A_exc_trap_inst_pri15_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_exc_trap_inst_pri15~q ),
	.prn(vcc));
defparam A_exc_trap_inst_pri15.is_wysiwyg = "true";
defparam A_exc_trap_inst_pri15.power_up = "low";

cyclonev_lcell_comb \A_exc_illegal_inst_pri15_nxt~0 (
	.dataa(!\M_exc_illegal_inst_pri15~q ),
	.datab(!\M_norm_intr_req~q ),
	.datac(!\hbreak_req~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_exc_illegal_inst_pri15_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_exc_illegal_inst_pri15_nxt~0 .extended_lut = "off";
defparam \A_exc_illegal_inst_pri15_nxt~0 .lut_mask = 64'hFDFDFDFDFDFDFDFD;
defparam \A_exc_illegal_inst_pri15_nxt~0 .shared_arith = "off";

dffeas A_exc_illegal_inst_pri15(
	.clk(clk_clk),
	.d(\A_exc_illegal_inst_pri15_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_exc_illegal_inst_pri15~q ),
	.prn(vcc));
defparam A_exc_illegal_inst_pri15.is_wysiwyg = "true";
defparam A_exc_illegal_inst_pri15.power_up = "low";

cyclonev_lcell_comb \A_exc_highest_pri_cause_code[0]~0 (
	.dataa(!\A_exc_norm_intr_pri5~q ),
	.datab(!\A_exc_trap_inst_pri15~q ),
	.datac(!\A_exc_illegal_inst_pri15~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_exc_highest_pri_cause_code[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_exc_highest_pri_cause_code[0]~0 .extended_lut = "off";
defparam \A_exc_highest_pri_cause_code[0]~0 .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \A_exc_highest_pri_cause_code[0]~0 .shared_arith = "off";

cyclonev_lcell_comb A_exc_active_no_break(
	.dataa(!\A_exc_any~q ),
	.datab(!\A_exc_allowed~q ),
	.datac(!\A_exc_break~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_exc_active_no_break~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam A_exc_active_no_break.extended_lut = "off";
defparam A_exc_active_no_break.lut_mask = 64'hF7F7F7F7F7F7F7F7;
defparam A_exc_active_no_break.shared_arith = "off";

dffeas \W_exception_reg_cause[0] (
	.clk(clk_clk),
	.d(\A_exc_highest_pri_cause_code[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_exc_active_no_break~combout ),
	.q(\W_exception_reg_cause[0]~q ),
	.prn(vcc));
defparam \W_exception_reg_cause[0] .is_wysiwyg = "true";
defparam \W_exception_reg_cause[0] .power_up = "low";

cyclonev_lcell_comb \E_control_reg_rddata_muxed[2]~2 (
	.dataa(!\Equal327~0_combout ),
	.datab(!\W_exception_reg_cause[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_control_reg_rddata_muxed[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_control_reg_rddata_muxed[2]~2 .extended_lut = "off";
defparam \E_control_reg_rddata_muxed[2]~2 .lut_mask = 64'h7777777777777777;
defparam \E_control_reg_rddata_muxed[2]~2 .shared_arith = "off";

dffeas \M_control_reg_rddata[2] (
	.clk(clk_clk),
	.d(\E_control_reg_rddata_muxed[2]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_control_reg_rddata[2]~q ),
	.prn(vcc));
defparam \M_control_reg_rddata[2] .is_wysiwyg = "true";
defparam \M_control_reg_rddata[2] .power_up = "low";

cyclonev_lcell_comb \M_inst_result[2]~2 (
	.dataa(!\M_exc_any~combout ),
	.datab(!\M_alu_result[2]~q ),
	.datac(!\M_ctrl_rd_ctl_reg~q ),
	.datad(!\M_pc_plus_one[0]~q ),
	.datae(!\M_control_reg_rddata[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_inst_result[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_inst_result[2]~2 .extended_lut = "off";
defparam \M_inst_result[2]~2 .lut_mask = 64'h7BFFFFFF7BFFFFFF;
defparam \M_inst_result[2]~2 .shared_arith = "off";

dffeas \A_inst_result[2] (
	.clk(clk_clk),
	.d(\M_inst_result[2]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_inst_result[2]~q ),
	.prn(vcc));
defparam \A_inst_result[2] .is_wysiwyg = "true";
defparam \A_inst_result[2] .power_up = "low";

dffeas \A_mul_cell_p1[2] (
	.clk(clk_clk),
	.d(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[2]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_mul_cell_p1[2]~q ),
	.prn(vcc));
defparam \A_mul_cell_p1[2] .is_wysiwyg = "true";
defparam \A_mul_cell_p1[2] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[2]~4 (
	.dataa(!\A_slow_inst_result[2]~q ),
	.datab(!\A_shift_rot_result[2]~q ),
	.datac(!\A_inst_result[2]~q ),
	.datad(!\A_mul_cell_p1[2]~q ),
	.datae(!\A_wr_data_unfiltered[15]~0_combout ),
	.dataf(!\A_wr_data_unfiltered[15]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[2]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[2]~4 .extended_lut = "off";
defparam \A_wr_data_unfiltered[2]~4 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_wr_data_unfiltered[2]~4 .shared_arith = "off";

dffeas \W_wr_data[2] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[2]~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[2]~q ),
	.prn(vcc));
defparam \W_wr_data[2] .is_wysiwyg = "true";
defparam \W_wr_data[2] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[2]~6 (
	.dataa(!\M_alu_result[2]~q ),
	.datab(!\A_wr_data_unfiltered[2]~4_combout ),
	.datac(!\first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[2] ),
	.datad(!\W_wr_data[2]~q ),
	.datae(!\E_src1[26]~0_combout ),
	.dataf(!\E_src1[26]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[2]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[2]~6 .extended_lut = "off";
defparam \D_src1_reg[2]~6 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[2]~6 .shared_arith = "off";

dffeas \E_src1[2] (
	.clk(clk_clk),
	.d(\D_src1_reg[2]~6_combout ),
	.asdata(\E_alu_result[2]~combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\Equal303~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(!\A_mem_stall~q ),
	.q(\E_src1[2]~q ),
	.prn(vcc));
defparam \E_src1[2] .is_wysiwyg = "true";
defparam \E_src1[2] .power_up = "low";

cyclonev_lcell_comb \E_alu_result~2 (
	.dataa(!\E_src2[2]~q ),
	.datab(!\E_src1[2]~q ),
	.datac(!\E_logic_op[1]~q ),
	.datad(!\E_logic_op[0]~q ),
	.datae(!\E_ctrl_logic~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result~2 .extended_lut = "off";
defparam \E_alu_result~2 .lut_mask = 64'h6996FFFF6996FFFF;
defparam \E_alu_result~2 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[2] (
	.dataa(!\Add9~57_sumout ),
	.datab(!\E_ctrl_retaddr~q ),
	.datac(!\E_alu_result~0_combout ),
	.datad(!\E_alu_result~2_combout ),
	.datae(!\E_extra_pc[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[2]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[2] .extended_lut = "off";
defparam \E_alu_result[2] .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \E_alu_result[2] .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[2]~14 (
	.dataa(!\D_src2_reg[0]~7_combout ),
	.datab(!\D_src2_reg[0]~8_combout ),
	.datac(!\W_wr_data[2]~q ),
	.datad(!\A_wr_data_unfiltered[2]~4_combout ),
	.datae(!\M_alu_result[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[2]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[2]~14 .extended_lut = "off";
defparam \D_src2_reg[2]~14 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \D_src2_reg[2]~14 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[2]~46 (
	.dataa(!\D_ctrl_src2_choose_imm~q ),
	.datab(!\E_src2[1]~0_combout ),
	.datac(!\D_iw[8]~q ),
	.datad(!\D_src2_reg[0]~4_combout ),
	.datae(!\D_src2_reg[2]~14_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[2]~46_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[2]~46 .extended_lut = "off";
defparam \D_src2[2]~46 .lut_mask = 64'h8DFFFFFF8DFFFFFF;
defparam \D_src2[2]~46 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[2]~8 (
	.dataa(!\D_ctrl_src2_choose_imm~q ),
	.datab(!\D_src2_reg[0]~4_combout ),
	.datac(!\D_src2_reg[0]~5_combout ),
	.datad(!\E_alu_result[2]~combout ),
	.datae(!\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[2] ),
	.dataf(!\D_src2[2]~46_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[2]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[2]~8 .extended_lut = "off";
defparam \D_src2[2]~8 .lut_mask = 64'h7DFFFFFFFFFFFFFF;
defparam \D_src2[2]~8 .shared_arith = "off";

dffeas \E_src2[2] (
	.clk(clk_clk),
	.d(\D_src2[2]~8_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_src2[2]~q ),
	.prn(vcc));
defparam \E_src2[2] .is_wysiwyg = "true";
defparam \E_src2[2] .power_up = "low";

cyclonev_lcell_comb \E_rot_mask[4]~4 (
	.dataa(!\E_src2[2]~q ),
	.datab(!\E_src2[1]~q ),
	.datac(!\E_src2[0]~q ),
	.datad(!\E_ctrl_shift_rot_right~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_mask[4]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_mask[4]~4 .extended_lut = "off";
defparam \E_rot_mask[4]~4 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \E_rot_mask[4]~4 .shared_arith = "off";

dffeas \M_rot_mask[4] (
	.clk(clk_clk),
	.d(\E_rot_mask[4]~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_rot_mask[4]~q ),
	.prn(vcc));
defparam \M_rot_mask[4] .is_wysiwyg = "true";
defparam \M_rot_mask[4] .power_up = "low";

cyclonev_lcell_comb \M_rot[4]~4 (
	.dataa(!\M_rot_prestep2[4]~q ),
	.datab(!\M_rot_prestep2[28]~q ),
	.datac(!\M_rot_prestep2[20]~q ),
	.datad(!\M_rot_prestep2[12]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[4]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[4]~4 .extended_lut = "off";
defparam \M_rot[4]~4 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[4]~4 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~4 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_pass0~q ),
	.datac(!\M_rot_sel_fill0~q ),
	.datad(!\M_rot_mask[4]~q ),
	.datae(!\M_rot[4]~4_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~4 .extended_lut = "off";
defparam \A_shift_rot_result~4 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~4 .shared_arith = "off";

dffeas \A_shift_rot_result[4] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_shift_rot_result[4]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[4] .is_wysiwyg = "true";
defparam \A_shift_rot_result[4] .power_up = "low";

cyclonev_lcell_comb \A_exc_highest_pri_cause_code[1]~1 (
	.dataa(!\A_exc_norm_intr_pri5~q ),
	.datab(!\A_exc_trap_inst_pri15~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_exc_highest_pri_cause_code[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_exc_highest_pri_cause_code[1]~1 .extended_lut = "off";
defparam \A_exc_highest_pri_cause_code[1]~1 .lut_mask = 64'h7777777777777777;
defparam \A_exc_highest_pri_cause_code[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \W_exception_reg_cause[2]~0 (
	.dataa(!\A_exc_highest_pri_cause_code[1]~1_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_exception_reg_cause[2]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_exception_reg_cause[2]~0 .extended_lut = "off";
defparam \W_exception_reg_cause[2]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \W_exception_reg_cause[2]~0 .shared_arith = "off";

dffeas \W_exception_reg_cause[2] (
	.clk(clk_clk),
	.d(\W_exception_reg_cause[2]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_exc_active_no_break~combout ),
	.q(\W_exception_reg_cause[2]~q ),
	.prn(vcc));
defparam \W_exception_reg_cause[2] .is_wysiwyg = "true";
defparam \W_exception_reg_cause[2] .power_up = "low";

cyclonev_lcell_comb \E_control_reg_rddata_muxed[4]~4 (
	.dataa(!\Equal327~0_combout ),
	.datab(!\W_exception_reg_cause[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_control_reg_rddata_muxed[4]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_control_reg_rddata_muxed[4]~4 .extended_lut = "off";
defparam \E_control_reg_rddata_muxed[4]~4 .lut_mask = 64'h7777777777777777;
defparam \E_control_reg_rddata_muxed[4]~4 .shared_arith = "off";

dffeas \M_control_reg_rddata[4] (
	.clk(clk_clk),
	.d(\E_control_reg_rddata_muxed[4]~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_control_reg_rddata[4]~q ),
	.prn(vcc));
defparam \M_control_reg_rddata[4] .is_wysiwyg = "true";
defparam \M_control_reg_rddata[4] .power_up = "low";

cyclonev_lcell_comb \M_inst_result[4]~4 (
	.dataa(!\M_exc_any~combout ),
	.datab(!\M_alu_result[4]~q ),
	.datac(!\M_ctrl_rd_ctl_reg~q ),
	.datad(!\M_pc_plus_one[2]~q ),
	.datae(!\M_control_reg_rddata[4]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_inst_result[4]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_inst_result[4]~4 .extended_lut = "off";
defparam \M_inst_result[4]~4 .lut_mask = 64'h7BFFFFFF7BFFFFFF;
defparam \M_inst_result[4]~4 .shared_arith = "off";

dffeas \A_inst_result[4] (
	.clk(clk_clk),
	.d(\M_inst_result[4]~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_inst_result[4]~q ),
	.prn(vcc));
defparam \A_inst_result[4] .is_wysiwyg = "true";
defparam \A_inst_result[4] .power_up = "low";

dffeas \A_mul_cell_p1[4] (
	.clk(clk_clk),
	.d(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[4]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_mul_cell_p1[4]~q ),
	.prn(vcc));
defparam \A_mul_cell_p1[4] .is_wysiwyg = "true";
defparam \A_mul_cell_p1[4] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[4]~6 (
	.dataa(!\A_slow_inst_result[4]~q ),
	.datab(!\A_shift_rot_result[4]~q ),
	.datac(!\A_inst_result[4]~q ),
	.datad(!\A_mul_cell_p1[4]~q ),
	.datae(!\A_wr_data_unfiltered[15]~0_combout ),
	.dataf(!\A_wr_data_unfiltered[15]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[4]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[4]~6 .extended_lut = "off";
defparam \A_wr_data_unfiltered[4]~6 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_wr_data_unfiltered[4]~6 .shared_arith = "off";

dffeas \W_wr_data[4] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[4]~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[4]~q ),
	.prn(vcc));
defparam \W_wr_data[4] .is_wysiwyg = "true";
defparam \W_wr_data[4] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[4]~16 (
	.dataa(!\M_alu_result[4]~q ),
	.datab(!\A_wr_data_unfiltered[4]~6_combout ),
	.datac(!\first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[4] ),
	.datad(!\W_wr_data[4]~q ),
	.datae(!\E_src1[26]~0_combout ),
	.dataf(!\E_src1[26]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[4]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[4]~16 .extended_lut = "off";
defparam \D_src1_reg[4]~16 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[4]~16 .shared_arith = "off";

dffeas \E_src1[4] (
	.clk(clk_clk),
	.d(\D_src1_reg[4]~16_combout ),
	.asdata(\E_alu_result[4]~combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\Equal303~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(!\A_mem_stall~q ),
	.q(\E_src1[4]~q ),
	.prn(vcc));
defparam \E_src1[4] .is_wysiwyg = "true";
defparam \E_src1[4] .power_up = "low";

cyclonev_lcell_comb \E_alu_result~3 (
	.dataa(!\E_src2[4]~q ),
	.datab(!\E_src1[4]~q ),
	.datac(!\E_logic_op[1]~q ),
	.datad(!\E_logic_op[0]~q ),
	.datae(!\E_ctrl_logic~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result~3 .extended_lut = "off";
defparam \E_alu_result~3 .lut_mask = 64'h6996FFFF6996FFFF;
defparam \E_alu_result~3 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[4] (
	.dataa(!\Add9~1_sumout ),
	.datab(!\E_ctrl_retaddr~q ),
	.datac(!\E_alu_result~0_combout ),
	.datad(!\E_alu_result~3_combout ),
	.datae(!\E_extra_pc[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[4]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[4] .extended_lut = "off";
defparam \E_alu_result[4] .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \E_alu_result[4] .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[4]~18 (
	.dataa(!\D_src2_reg[0]~7_combout ),
	.datab(!\D_src2_reg[0]~8_combout ),
	.datac(!\W_wr_data[4]~q ),
	.datad(!\A_wr_data_unfiltered[4]~6_combout ),
	.datae(!\M_alu_result[4]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[4]~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[4]~18 .extended_lut = "off";
defparam \D_src2_reg[4]~18 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \D_src2_reg[4]~18 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[4]~43 (
	.dataa(!\D_ctrl_src2_choose_imm~q ),
	.datab(!\E_src2[1]~0_combout ),
	.datac(!\D_iw[10]~q ),
	.datad(!\D_src2_reg[0]~4_combout ),
	.datae(!\D_src2_reg[4]~18_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[4]~43_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[4]~43 .extended_lut = "off";
defparam \D_src2[4]~43 .lut_mask = 64'h8DFFFFFF8DFFFFFF;
defparam \D_src2[4]~43 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[4]~16 (
	.dataa(!\D_ctrl_src2_choose_imm~q ),
	.datab(!\D_src2_reg[0]~4_combout ),
	.datac(!\D_src2_reg[0]~5_combout ),
	.datad(!\E_alu_result[4]~combout ),
	.datae(!\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[4] ),
	.dataf(!\D_src2[4]~43_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[4]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[4]~16 .extended_lut = "off";
defparam \D_src2[4]~16 .lut_mask = 64'h7DFFFFFFFFFFFFFF;
defparam \D_src2[4]~16 .shared_arith = "off";

dffeas \E_src2[4] (
	.clk(clk_clk),
	.d(\D_src2[4]~16_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_src2[4]~q ),
	.prn(vcc));
defparam \E_src2[4] .is_wysiwyg = "true";
defparam \E_src2[4] .power_up = "low";

cyclonev_lcell_comb \E_rot_sel_fill0~0 (
	.dataa(!\E_src2[3]~q ),
	.datab(!\E_src2[4]~q ),
	.datac(!\E_ctrl_shift_rot_left~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_sel_fill0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_sel_fill0~0 .extended_lut = "off";
defparam \E_rot_sel_fill0~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \E_rot_sel_fill0~0 .shared_arith = "off";

dffeas M_rot_sel_fill0(
	.clk(clk_clk),
	.d(\E_rot_sel_fill0~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_rot_sel_fill0~q ),
	.prn(vcc));
defparam M_rot_sel_fill0.is_wysiwyg = "true";
defparam M_rot_sel_fill0.power_up = "low";

cyclonev_lcell_comb \M_rot[3]~3 (
	.dataa(!\M_rot_prestep2[3]~q ),
	.datab(!\M_rot_prestep2[27]~q ),
	.datac(!\M_rot_prestep2[19]~q ),
	.datad(!\M_rot_prestep2[11]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[3]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[3]~3 .extended_lut = "off";
defparam \M_rot[3]~3 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[3]~3 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~3 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_pass0~q ),
	.datac(!\M_rot_sel_fill0~q ),
	.datad(!\M_rot_mask[3]~q ),
	.datae(!\M_rot[3]~3_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~3 .extended_lut = "off";
defparam \A_shift_rot_result~3 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~3 .shared_arith = "off";

dffeas \A_shift_rot_result[3] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_shift_rot_result[3]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[3] .is_wysiwyg = "true";
defparam \A_shift_rot_result[3] .power_up = "low";

dffeas \W_exception_reg_cause[1] (
	.clk(clk_clk),
	.d(\A_exc_highest_pri_cause_code[1]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_exc_active_no_break~combout ),
	.q(\W_exception_reg_cause[1]~q ),
	.prn(vcc));
defparam \W_exception_reg_cause[1] .is_wysiwyg = "true";
defparam \W_exception_reg_cause[1] .power_up = "low";

cyclonev_lcell_comb \E_control_reg_rddata_muxed[3]~3 (
	.dataa(!\Equal327~0_combout ),
	.datab(!\W_exception_reg_cause[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_control_reg_rddata_muxed[3]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_control_reg_rddata_muxed[3]~3 .extended_lut = "off";
defparam \E_control_reg_rddata_muxed[3]~3 .lut_mask = 64'h7777777777777777;
defparam \E_control_reg_rddata_muxed[3]~3 .shared_arith = "off";

dffeas \M_control_reg_rddata[3] (
	.clk(clk_clk),
	.d(\E_control_reg_rddata_muxed[3]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_control_reg_rddata[3]~q ),
	.prn(vcc));
defparam \M_control_reg_rddata[3] .is_wysiwyg = "true";
defparam \M_control_reg_rddata[3] .power_up = "low";

cyclonev_lcell_comb \M_inst_result[3]~3 (
	.dataa(!\M_exc_any~combout ),
	.datab(!\M_alu_result[3]~q ),
	.datac(!\M_ctrl_rd_ctl_reg~q ),
	.datad(!\M_pc_plus_one[1]~q ),
	.datae(!\M_control_reg_rddata[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_inst_result[3]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_inst_result[3]~3 .extended_lut = "off";
defparam \M_inst_result[3]~3 .lut_mask = 64'h7BFFFFFF7BFFFFFF;
defparam \M_inst_result[3]~3 .shared_arith = "off";

dffeas \A_inst_result[3] (
	.clk(clk_clk),
	.d(\M_inst_result[3]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_inst_result[3]~q ),
	.prn(vcc));
defparam \A_inst_result[3] .is_wysiwyg = "true";
defparam \A_inst_result[3] .power_up = "low";

dffeas \A_mul_cell_p1[3] (
	.clk(clk_clk),
	.d(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[3]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_mul_cell_p1[3]~q ),
	.prn(vcc));
defparam \A_mul_cell_p1[3] .is_wysiwyg = "true";
defparam \A_mul_cell_p1[3] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[3]~5 (
	.dataa(!\A_slow_inst_result[3]~q ),
	.datab(!\A_shift_rot_result[3]~q ),
	.datac(!\A_inst_result[3]~q ),
	.datad(!\A_mul_cell_p1[3]~q ),
	.datae(!\A_wr_data_unfiltered[15]~0_combout ),
	.dataf(!\A_wr_data_unfiltered[15]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[3]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[3]~5 .extended_lut = "off";
defparam \A_wr_data_unfiltered[3]~5 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_wr_data_unfiltered[3]~5 .shared_arith = "off";

dffeas \W_wr_data[3] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[3]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[3]~q ),
	.prn(vcc));
defparam \W_wr_data[3] .is_wysiwyg = "true";
defparam \W_wr_data[3] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[3]~0 (
	.dataa(!\M_alu_result[3]~q ),
	.datab(!\A_wr_data_unfiltered[3]~5_combout ),
	.datac(!\first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[3] ),
	.datad(!\W_wr_data[3]~q ),
	.datae(!\E_src1[26]~0_combout ),
	.dataf(!\E_src1[26]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[3]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[3]~0 .extended_lut = "off";
defparam \D_src1_reg[3]~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[3]~0 .shared_arith = "off";

dffeas \E_src1[3] (
	.clk(clk_clk),
	.d(\D_src1_reg[3]~0_combout ),
	.asdata(\E_alu_result[3]~combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\Equal303~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(!\A_mem_stall~q ),
	.q(\E_src1[3]~q ),
	.prn(vcc));
defparam \E_src1[3] .is_wysiwyg = "true";
defparam \E_src1[3] .power_up = "low";

cyclonev_lcell_comb \E_alu_result[3] (
	.dataa(!\Add9~53_sumout ),
	.datab(!\E_ctrl_cmp~q ),
	.datac(!\E_logic_result[3]~0_combout ),
	.datad(!\E_ctrl_logic~q ),
	.datae(!\E_ctrl_retaddr~q ),
	.dataf(!\E_extra_pc[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[3]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[3] .extended_lut = "off";
defparam \E_alu_result[3] .lut_mask = 64'hDFFFFFDFFFFFFFFF;
defparam \E_alu_result[3] .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[3]~16 (
	.dataa(!\D_src2_reg[0]~7_combout ),
	.datab(!\D_src2_reg[0]~8_combout ),
	.datac(!\W_wr_data[3]~q ),
	.datad(!\A_wr_data_unfiltered[3]~5_combout ),
	.datae(!\M_alu_result[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[3]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[3]~16 .extended_lut = "off";
defparam \D_src2_reg[3]~16 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \D_src2_reg[3]~16 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[3]~45 (
	.dataa(!\D_ctrl_src2_choose_imm~q ),
	.datab(!\E_src2[1]~0_combout ),
	.datac(!\D_iw[9]~q ),
	.datad(!\D_src2_reg[0]~4_combout ),
	.datae(!\D_src2_reg[3]~16_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[3]~45_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[3]~45 .extended_lut = "off";
defparam \D_src2[3]~45 .lut_mask = 64'h8DFFFFFF8DFFFFFF;
defparam \D_src2[3]~45 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[3]~0 (
	.dataa(!\D_ctrl_src2_choose_imm~q ),
	.datab(!\D_src2_reg[0]~4_combout ),
	.datac(!\D_src2_reg[0]~5_combout ),
	.datad(!\E_alu_result[3]~combout ),
	.datae(!\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[3] ),
	.dataf(!\D_src2[3]~45_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[3]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[3]~0 .extended_lut = "off";
defparam \D_src2[3]~0 .lut_mask = 64'h7DFFFFFFFFFFFFFF;
defparam \D_src2[3]~0 .shared_arith = "off";

dffeas \E_src2[3] (
	.clk(clk_clk),
	.d(\D_src2[3]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_src2[3]~q ),
	.prn(vcc));
defparam \E_src2[3] .is_wysiwyg = "true";
defparam \E_src2[3] .power_up = "low";

cyclonev_lcell_comb \E_rot_pass0~0 (
	.dataa(!\E_src2[3]~q ),
	.datab(!\E_src2[4]~q ),
	.datac(!\E_ctrl_rot~q ),
	.datad(!\E_ctrl_shift_rot_right~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_pass0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_pass0~0 .extended_lut = "off";
defparam \E_rot_pass0~0 .lut_mask = 64'hEFFFEFFFEFFFEFFF;
defparam \E_rot_pass0~0 .shared_arith = "off";

dffeas M_rot_pass0(
	.clk(clk_clk),
	.d(\E_rot_pass0~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_rot_pass0~q ),
	.prn(vcc));
defparam M_rot_pass0.is_wysiwyg = "true";
defparam M_rot_pass0.power_up = "low";

cyclonev_lcell_comb \M_rot[0]~0 (
	.dataa(!\M_rot_prestep2[0]~q ),
	.datab(!\M_rot_prestep2[24]~q ),
	.datac(!\M_rot_prestep2[16]~q ),
	.datad(!\M_rot_prestep2[8]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[0]~0 .extended_lut = "off";
defparam \M_rot[0]~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~0 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_pass0~q ),
	.datac(!\M_rot_mask[0]~q ),
	.datad(!\M_rot_sel_fill0~q ),
	.datae(!\M_rot[0]~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~0 .extended_lut = "off";
defparam \A_shift_rot_result~0 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~0 .shared_arith = "off";

dffeas \A_shift_rot_result[0] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_shift_rot_result[0]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[0] .is_wysiwyg = "true";
defparam \A_shift_rot_result[0] .power_up = "low";

cyclonev_lcell_comb \W_estatus_reg_pie_nxt~0 (
	.dataa(!\A_valid_from_M~q ),
	.datab(!\A_iw[7]~q ),
	.datac(!\A_iw[6]~q ),
	.datad(!\A_wrctl_status~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_estatus_reg_pie_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_estatus_reg_pie_nxt~0 .extended_lut = "off";
defparam \W_estatus_reg_pie_nxt~0 .lut_mask = 64'hDFFFDFFFDFFFDFFF;
defparam \W_estatus_reg_pie_nxt~0 .shared_arith = "off";

cyclonev_lcell_comb \W_estatus_reg_pie_nxt~1 (
	.dataa(!\W_status_reg_pie~q ),
	.datab(!\A_inst_result[0]~q ),
	.datac(!\W_estatus_reg_pie~q ),
	.datad(!\A_exc_active_no_break~combout ),
	.datae(!\W_estatus_reg_pie_nxt~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_estatus_reg_pie_nxt~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_estatus_reg_pie_nxt~1 .extended_lut = "off";
defparam \W_estatus_reg_pie_nxt~1 .lut_mask = 64'h7FFFFF7F7FFFFF7F;
defparam \W_estatus_reg_pie_nxt~1 .shared_arith = "off";

dffeas W_estatus_reg_pie(
	.clk(clk_clk),
	.d(\W_estatus_reg_pie_nxt~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_estatus_reg_pie~q ),
	.prn(vcc));
defparam W_estatus_reg_pie.is_wysiwyg = "true";
defparam W_estatus_reg_pie.power_up = "low";

cyclonev_lcell_comb \W_bstatus_reg_pie_nxt~0 (
	.dataa(!\A_valid_from_M~q ),
	.datab(!\A_iw[7]~q ),
	.datac(!\A_iw[6]~q ),
	.datad(!\A_wrctl_status~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_bstatus_reg_pie_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_bstatus_reg_pie_nxt~0 .extended_lut = "off";
defparam \W_bstatus_reg_pie_nxt~0 .lut_mask = 64'hF7FFF7FFF7FFF7FF;
defparam \W_bstatus_reg_pie_nxt~0 .shared_arith = "off";

cyclonev_lcell_comb \W_bstatus_reg_pie_nxt~1 (
	.dataa(!\A_exc_allowed~q ),
	.datab(!\W_status_reg_pie~q ),
	.datac(!\A_exc_break~q ),
	.datad(!\A_inst_result[0]~q ),
	.datae(!\W_bstatus_reg_pie~q ),
	.dataf(!\W_bstatus_reg_pie_nxt~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_bstatus_reg_pie_nxt~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_bstatus_reg_pie_nxt~1 .extended_lut = "off";
defparam \W_bstatus_reg_pie_nxt~1 .lut_mask = 64'hB7FFFFFF7BFFFFFF;
defparam \W_bstatus_reg_pie_nxt~1 .shared_arith = "off";

dffeas W_bstatus_reg_pie(
	.clk(clk_clk),
	.d(\W_bstatus_reg_pie_nxt~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_bstatus_reg_pie~q ),
	.prn(vcc));
defparam W_bstatus_reg_pie.is_wysiwyg = "true";
defparam W_bstatus_reg_pie.power_up = "low";

cyclonev_lcell_comb \D_control_reg_rddata_muxed[0]~0 (
	.dataa(!\W_status_reg_pie~q ),
	.datab(!\W_estatus_reg_pie~q ),
	.datac(!\W_bstatus_reg_pie~q ),
	.datad(!\D_iw[6]~q ),
	.datae(!\D_iw[7]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_control_reg_rddata_muxed[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_control_reg_rddata_muxed[0]~0 .extended_lut = "off";
defparam \D_control_reg_rddata_muxed[0]~0 .lut_mask = 64'h7FFFFF7F7FFFFF7F;
defparam \D_control_reg_rddata_muxed[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \D_control_reg_rddata_muxed[0]~1 (
	.dataa(!\D_iw[10]~q ),
	.datab(!\D_iw[8]~q ),
	.datac(!\D_iw[9]~q ),
	.datad(!\D_control_reg_rddata_muxed[0]~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_control_reg_rddata_muxed[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_control_reg_rddata_muxed[0]~1 .extended_lut = "off";
defparam \D_control_reg_rddata_muxed[0]~1 .lut_mask = 64'hFEFFFEFFFEFFFEFF;
defparam \D_control_reg_rddata_muxed[0]~1 .shared_arith = "off";

dffeas \E_control_reg_rddata[0] (
	.clk(clk_clk),
	.d(\D_control_reg_rddata_muxed[0]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_control_reg_rddata[0]~q ),
	.prn(vcc));
defparam \E_control_reg_rddata[0] .is_wysiwyg = "true";
defparam \E_control_reg_rddata[0] .power_up = "low";

cyclonev_lcell_comb \E_control_reg_rddata_muxed[0]~0 (
	.dataa(!\E_control_reg_rddata[0]~q ),
	.datab(!\M_control_reg_rddata[16]~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_control_reg_rddata_muxed[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_control_reg_rddata_muxed[0]~0 .extended_lut = "off";
defparam \E_control_reg_rddata_muxed[0]~0 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \E_control_reg_rddata_muxed[0]~0 .shared_arith = "off";

dffeas \M_control_reg_rddata[0] (
	.clk(clk_clk),
	.d(\E_control_reg_rddata_muxed[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_control_reg_rddata[0]~q ),
	.prn(vcc));
defparam \M_control_reg_rddata[0] .is_wysiwyg = "true";
defparam \M_control_reg_rddata[0] .power_up = "low";

cyclonev_lcell_comb \M_inst_result[0]~0 (
	.dataa(!\M_exc_any~combout ),
	.datab(!\M_alu_result[0]~q ),
	.datac(!\M_control_reg_rddata[0]~q ),
	.datad(!\M_ctrl_rd_ctl_reg~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_inst_result[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_inst_result[0]~0 .extended_lut = "off";
defparam \M_inst_result[0]~0 .lut_mask = 64'hAF3FAF3FAF3FAF3F;
defparam \M_inst_result[0]~0 .shared_arith = "off";

dffeas \A_inst_result[0] (
	.clk(clk_clk),
	.d(\M_inst_result[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_inst_result[0]~q ),
	.prn(vcc));
defparam \A_inst_result[0] .is_wysiwyg = "true";
defparam \A_inst_result[0] .power_up = "low";

dffeas \A_mul_cell_p1[0] (
	.clk(clk_clk),
	.d(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[0]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_mul_cell_p1[0]~q ),
	.prn(vcc));
defparam \A_mul_cell_p1[0] .is_wysiwyg = "true";
defparam \A_mul_cell_p1[0] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[0]~2 (
	.dataa(!\A_slow_inst_result[0]~q ),
	.datab(!\A_shift_rot_result[0]~q ),
	.datac(!\A_inst_result[0]~q ),
	.datad(!\A_mul_cell_p1[0]~q ),
	.datae(!\A_wr_data_unfiltered[15]~0_combout ),
	.dataf(!\A_wr_data_unfiltered[15]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[0]~2 .extended_lut = "off";
defparam \A_wr_data_unfiltered[0]~2 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_wr_data_unfiltered[0]~2 .shared_arith = "off";

dffeas \W_wr_data[0] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[0]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[0]~q ),
	.prn(vcc));
defparam \W_wr_data[0] .is_wysiwyg = "true";
defparam \W_wr_data[0] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[0]~10 (
	.dataa(!\W_wr_data[0]~q ),
	.datab(!\D_src2_reg[0]~7_combout ),
	.datac(!\A_wr_data_unfiltered[0]~2_combout ),
	.datad(!\D_src2_reg[0]~8_combout ),
	.datae(!\M_alu_result[0]~q ),
	.dataf(!\D_src2_reg[0]~9_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[0]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[0]~10 .extended_lut = "off";
defparam \D_src2_reg[0]~10 .lut_mask = 64'h7FDFFFFFFFFFFFFF;
defparam \D_src2_reg[0]~10 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[0]~47 (
	.dataa(!\E_src2[1]~0_combout ),
	.datab(!\D_src2_reg[0]~6_combout ),
	.datac(!\D_iw[6]~q ),
	.datad(!\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[0] ),
	.datae(!\D_ctrl_src2_choose_imm~q ),
	.dataf(!\D_src2_reg[0]~3_combout ),
	.datag(!\D_src2_reg[0]~10_combout ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[0]~47_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[0]~47 .extended_lut = "on";
defparam \D_src2[0]~47 .lut_mask = 64'hFFFDFFFDFFFDFFFD;
defparam \D_src2[0]~47 .shared_arith = "off";

dffeas \E_src2[0] (
	.clk(clk_clk),
	.d(\D_src2[0]~47_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_src2[0]~q ),
	.prn(vcc));
defparam \E_src2[0] .is_wysiwyg = "true";
defparam \E_src2[0] .power_up = "low";

dffeas \M_mem_baddr[0] (
	.clk(clk_clk),
	.d(\Add9~65_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_mem_baddr[0]~q ),
	.prn(vcc));
defparam \M_mem_baddr[0] .is_wysiwyg = "true";
defparam \M_mem_baddr[0] .power_up = "low";

cyclonev_lcell_comb M_ld_align_sh8(
	.dataa(!\M_mem_baddr[0]~q ),
	.datab(!\M_ld_align_byte1_fill~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_ld_align_sh8~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam M_ld_align_sh8.extended_lut = "off";
defparam M_ld_align_sh8.lut_mask = 64'h7777777777777777;
defparam M_ld_align_sh8.shared_arith = "off";

dffeas A_ld_align_sh8(
	.clk(clk_clk),
	.d(\M_ld_align_sh8~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_ld_align_sh8~q ),
	.prn(vcc));
defparam A_ld_align_sh8.is_wysiwyg = "true";
defparam A_ld_align_sh8.power_up = "low";

cyclonev_lcell_comb \A_slow_inst_result_nxt[1]~1 (
	.dataa(!\d_readdata_d1[1]~q ),
	.datab(!\d_readdata_d1[17]~q ),
	.datac(!\d_readdata_d1[9]~q ),
	.datad(!\d_readdata_d1[25]~q ),
	.datae(!\A_ld_align_sh16~q ),
	.dataf(!\A_ld_align_sh8~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[1]~1 .extended_lut = "off";
defparam \A_slow_inst_result_nxt[1]~1 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_slow_inst_result_nxt[1]~1 .shared_arith = "off";

dffeas \A_slow_inst_result[1] (
	.clk(clk_clk),
	.d(\A_slow_inst_result_nxt[1]~1_combout ),
	.asdata(d_readdata[1]),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_ctrl_ld32~q ),
	.ena(\A_ctrl_ld~q ),
	.q(\A_slow_inst_result[1]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[1] .is_wysiwyg = "true";
defparam \A_slow_inst_result[1] .power_up = "low";

cyclonev_lcell_comb \M_rot[1]~1 (
	.dataa(!\M_rot_prestep2[1]~q ),
	.datab(!\M_rot_prestep2[25]~q ),
	.datac(!\M_rot_prestep2[17]~q ),
	.datad(!\M_rot_prestep2[9]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[1]~1 .extended_lut = "off";
defparam \M_rot[1]~1 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~1 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_pass0~q ),
	.datac(!\M_rot_sel_fill0~q ),
	.datad(!\M_rot_mask[1]~q ),
	.datae(!\M_rot[1]~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~1 .extended_lut = "off";
defparam \A_shift_rot_result~1 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~1 .shared_arith = "off";

dffeas \A_shift_rot_result[1] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_shift_rot_result[1]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[1] .is_wysiwyg = "true";
defparam \A_shift_rot_result[1] .power_up = "low";

dffeas W_ienable_reg_irq1(
	.clk(clk_clk),
	.d(\A_inst_result[1]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_ienable_reg_irq1_nxt~0_combout ),
	.q(\W_ienable_reg_irq1~q ),
	.prn(vcc));
defparam W_ienable_reg_irq1.is_wysiwyg = "true";
defparam W_ienable_reg_irq1.power_up = "low";

cyclonev_lcell_comb W_ipending_reg_irq1_nxt(
	.dataa(!\W_ienable_reg_irq1~q ),
	.datab(!\the_first_nios2_system_cpu_cpu_nios2_oci|the_first_nios2_system_cpu_cpu_nios2_avalon_reg|oci_ienable[1]~q ),
	.datac(!timeout_occurred),
	.datad(!control_register_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_ipending_reg_irq1_nxt~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam W_ipending_reg_irq1_nxt.extended_lut = "off";
defparam W_ipending_reg_irq1_nxt.lut_mask = 64'hDFFFDFFFDFFFDFFF;
defparam W_ipending_reg_irq1_nxt.shared_arith = "off";

dffeas W_ipending_reg_irq1(
	.clk(clk_clk),
	.d(\W_ipending_reg_irq1_nxt~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_ipending_reg_irq1~q ),
	.prn(vcc));
defparam W_ipending_reg_irq1.is_wysiwyg = "true";
defparam W_ipending_reg_irq1.power_up = "low";

cyclonev_lcell_comb \D_control_reg_rddata_muxed[1]~2 (
	.dataa(!\W_ipending_reg_irq1~q ),
	.datab(!\W_ienable_reg_irq1~q ),
	.datac(!\Equal324~0_combout ),
	.datad(!\E_control_reg_rddata[1]~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_control_reg_rddata_muxed[1]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_control_reg_rddata_muxed[1]~2 .extended_lut = "off";
defparam \D_control_reg_rddata_muxed[1]~2 .lut_mask = 64'h53FF53FF53FF53FF;
defparam \D_control_reg_rddata_muxed[1]~2 .shared_arith = "off";

dffeas \E_control_reg_rddata[1] (
	.clk(clk_clk),
	.d(\D_control_reg_rddata_muxed[1]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_control_reg_rddata[1]~q ),
	.prn(vcc));
defparam \E_control_reg_rddata[1] .is_wysiwyg = "true";
defparam \E_control_reg_rddata[1] .power_up = "low";

cyclonev_lcell_comb \E_control_reg_rddata_muxed[1]~1 (
	.dataa(!\M_control_reg_rddata[16]~0_combout ),
	.datab(!\E_control_reg_rddata[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_control_reg_rddata_muxed[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_control_reg_rddata_muxed[1]~1 .extended_lut = "off";
defparam \E_control_reg_rddata_muxed[1]~1 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \E_control_reg_rddata_muxed[1]~1 .shared_arith = "off";

dffeas \M_control_reg_rddata[1] (
	.clk(clk_clk),
	.d(\E_control_reg_rddata_muxed[1]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_control_reg_rddata[1]~q ),
	.prn(vcc));
defparam \M_control_reg_rddata[1] .is_wysiwyg = "true";
defparam \M_control_reg_rddata[1] .power_up = "low";

cyclonev_lcell_comb \M_inst_result[1]~1 (
	.dataa(!\M_exc_any~combout ),
	.datab(!\M_alu_result[1]~q ),
	.datac(!\M_ctrl_rd_ctl_reg~q ),
	.datad(!\M_control_reg_rddata[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_inst_result[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_inst_result[1]~1 .extended_lut = "off";
defparam \M_inst_result[1]~1 .lut_mask = 64'hA3FFA3FFA3FFA3FF;
defparam \M_inst_result[1]~1 .shared_arith = "off";

dffeas \A_inst_result[1] (
	.clk(clk_clk),
	.d(\M_inst_result[1]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_inst_result[1]~q ),
	.prn(vcc));
defparam \A_inst_result[1] .is_wysiwyg = "true";
defparam \A_inst_result[1] .power_up = "low";

dffeas \A_mul_cell_p1[1] (
	.clk(clk_clk),
	.d(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[1]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_mul_cell_p1[1]~q ),
	.prn(vcc));
defparam \A_mul_cell_p1[1] .is_wysiwyg = "true";
defparam \A_mul_cell_p1[1] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[1]~3 (
	.dataa(!\A_slow_inst_result[1]~q ),
	.datab(!\A_shift_rot_result[1]~q ),
	.datac(!\A_inst_result[1]~q ),
	.datad(!\A_mul_cell_p1[1]~q ),
	.datae(!\A_wr_data_unfiltered[15]~0_combout ),
	.dataf(!\A_wr_data_unfiltered[15]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[1]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[1]~3 .extended_lut = "off";
defparam \A_wr_data_unfiltered[1]~3 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_wr_data_unfiltered[1]~3 .shared_arith = "off";

dffeas \W_wr_data[1] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[1]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[1]~q ),
	.prn(vcc));
defparam \W_wr_data[1] .is_wysiwyg = "true";
defparam \W_wr_data[1] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[1]~24 (
	.dataa(!\M_alu_result[1]~q ),
	.datab(!\A_wr_data_unfiltered[1]~3_combout ),
	.datac(!\first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[1] ),
	.datad(!\W_wr_data[1]~q ),
	.datae(!\E_src1[26]~0_combout ),
	.dataf(!\E_src1[26]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[1]~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[1]~24 .extended_lut = "off";
defparam \D_src1_reg[1]~24 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[1]~24 .shared_arith = "off";

dffeas \E_src1[1] (
	.clk(clk_clk),
	.d(\D_src1_reg[1]~24_combout ),
	.asdata(\E_alu_result[1]~combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\Equal303~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(!\A_mem_stall~q ),
	.q(\E_src1[1]~q ),
	.prn(vcc));
defparam \E_src1[1] .is_wysiwyg = "true";
defparam \E_src1[1] .power_up = "low";

cyclonev_lcell_comb \E_logic_result[1]~7 (
	.dataa(!\E_src2[1]~q ),
	.datab(!\E_src1[1]~q ),
	.datac(!\E_logic_op[1]~q ),
	.datad(!\E_logic_op[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[1]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[1]~7 .extended_lut = "off";
defparam \E_logic_result[1]~7 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[1]~7 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[1] (
	.dataa(!\E_logic_result[1]~7_combout ),
	.datab(!\E_ctrl_logic~q ),
	.datac(!\E_alu_result~0_combout ),
	.datad(!\Add9~69_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[1]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[1] .extended_lut = "off";
defparam \E_alu_result[1] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \E_alu_result[1] .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[1]~12 (
	.dataa(!\D_src2_reg[0]~7_combout ),
	.datab(!\D_src2_reg[0]~8_combout ),
	.datac(!\W_wr_data[1]~q ),
	.datad(!\A_wr_data_unfiltered[1]~3_combout ),
	.datae(!\M_alu_result[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[1]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[1]~12 .extended_lut = "off";
defparam \D_src2_reg[1]~12 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \D_src2_reg[1]~12 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[1]~44 (
	.dataa(!\D_ctrl_src2_choose_imm~q ),
	.datab(!\E_src2[1]~0_combout ),
	.datac(!\D_iw[7]~q ),
	.datad(!\D_src2_reg[0]~4_combout ),
	.datae(!\D_src2_reg[1]~12_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[1]~44_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[1]~44 .extended_lut = "off";
defparam \D_src2[1]~44 .lut_mask = 64'h8DFFFFFF8DFFFFFF;
defparam \D_src2[1]~44 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[1]~24 (
	.dataa(!\D_ctrl_src2_choose_imm~q ),
	.datab(!\D_src2_reg[0]~4_combout ),
	.datac(!\D_src2_reg[0]~5_combout ),
	.datad(!\E_alu_result[1]~combout ),
	.datae(!\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[1] ),
	.dataf(!\D_src2[1]~44_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[1]~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[1]~24 .extended_lut = "off";
defparam \D_src2[1]~24 .lut_mask = 64'h7DFFFFFFFFFFFFFF;
defparam \D_src2[1]~24 .shared_arith = "off";

dffeas \E_src2[1] (
	.clk(clk_clk),
	.d(\D_src2[1]~24_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_src2[1]~q ),
	.prn(vcc));
defparam \E_src2[1] .is_wysiwyg = "true";
defparam \E_src2[1] .power_up = "low";

dffeas \M_mem_baddr[1] (
	.clk(clk_clk),
	.d(\Add9~69_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_mem_baddr[1]~q ),
	.prn(vcc));
defparam \M_mem_baddr[1] .is_wysiwyg = "true";
defparam \M_mem_baddr[1] .power_up = "low";

dffeas \A_mem_baddr[1] (
	.clk(clk_clk),
	.d(\M_mem_baddr[1]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_mem_baddr[1]~q ),
	.prn(vcc));
defparam \A_mem_baddr[1] .is_wysiwyg = "true";
defparam \A_mem_baddr[1] .power_up = "low";

dffeas \A_mem_baddr[0] (
	.clk(clk_clk),
	.d(\M_mem_baddr[0]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_mem_baddr[0]~q ),
	.prn(vcc));
defparam \A_mem_baddr[0] .is_wysiwyg = "true";
defparam \A_mem_baddr[0] .power_up = "low";

dffeas A_ctrl_ld16(
	.clk(clk_clk),
	.d(\M_ctrl_ld16~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_ctrl_ld16~q ),
	.prn(vcc));
defparam A_ctrl_ld16.is_wysiwyg = "true";
defparam A_ctrl_ld16.power_up = "low";

cyclonev_lcell_comb \A_slow_ld_data_sign_bit~0 (
	.dataa(!\A_mem_baddr[0]~q ),
	.datab(!\A_ctrl_ld16~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_ld_data_sign_bit~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_ld_data_sign_bit~0 .extended_lut = "off";
defparam \A_slow_ld_data_sign_bit~0 .lut_mask = 64'h7777777777777777;
defparam \A_slow_ld_data_sign_bit~0 .shared_arith = "off";

dffeas M_ctrl_ld_signed(
	.clk(clk_clk),
	.d(\Equal219~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_ctrl_ld_signed~q ),
	.prn(vcc));
defparam M_ctrl_ld_signed.is_wysiwyg = "true";
defparam M_ctrl_ld_signed.power_up = "low";

dffeas A_ctrl_ld_signed(
	.clk(clk_clk),
	.d(\M_ctrl_ld_signed~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_ctrl_ld_signed~q ),
	.prn(vcc));
defparam A_ctrl_ld_signed.is_wysiwyg = "true";
defparam A_ctrl_ld_signed.power_up = "low";

cyclonev_lcell_comb \A_slow_ld_data_fill_bit~0 (
	.dataa(!\A_mem_baddr[1]~q ),
	.datab(!\d_readdata_d1[31]~q ),
	.datac(!\d_readdata_d1[15]~q ),
	.datad(!\d_readdata_d1[23]~q ),
	.datae(!\A_slow_ld_data_sign_bit~0_combout ),
	.dataf(!\A_ctrl_ld_signed~q ),
	.datag(!\d_readdata_d1[7]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_ld_data_fill_bit~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_ld_data_fill_bit~0 .extended_lut = "on";
defparam \A_slow_ld_data_fill_bit~0 .lut_mask = 64'hFFD8FFD8FFD8FFD8;
defparam \A_slow_ld_data_fill_bit~0 .shared_arith = "off";

cyclonev_lcell_comb \A_slow_inst_result_nxt[31]~38 (
	.dataa(!\A_ctrl_ld32~q ),
	.datab(!\A_ld_align_byte2_byte3_fill~q ),
	.datac(!src0_valid),
	.datad(!av_readdata_pre_31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[31]~38_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[31]~38 .extended_lut = "off";
defparam \A_slow_inst_result_nxt[31]~38 .lut_mask = 64'h27FF27FF27FF27FF;
defparam \A_slow_inst_result_nxt[31]~38 .shared_arith = "off";

cyclonev_lcell_comb \A_slow_inst_result_nxt[31]~12 (
	.dataa(!\A_ctrl_ld32~q ),
	.datab(!\d_readdata_d1[31]~q ),
	.datac(!\A_slow_ld_data_fill_bit~0_combout ),
	.datad(!src0_valid1),
	.datae(!q_a_31),
	.dataf(!\A_slow_inst_result_nxt[31]~38_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_nxt[31]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_nxt[31]~12 .extended_lut = "off";
defparam \A_slow_inst_result_nxt[31]~12 .lut_mask = 64'h7FFFFFFFBFFFFFFF;
defparam \A_slow_inst_result_nxt[31]~12 .shared_arith = "off";

dffeas \A_slow_inst_result[31] (
	.clk(clk_clk),
	.d(\A_slow_inst_result_nxt[31]~12_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_ctrl_ld~q ),
	.q(\A_slow_inst_result[31]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[31] .is_wysiwyg = "true";
defparam \A_slow_inst_result[31] .power_up = "low";

cyclonev_lcell_comb \M_rot[7]~12 (
	.dataa(!\M_rot_prestep2[31]~q ),
	.datab(!\M_rot_prestep2[23]~q ),
	.datac(!\M_rot_prestep2[15]~q ),
	.datad(!\M_rot_prestep2[7]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[7]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[7]~12 .extended_lut = "off";
defparam \M_rot[7]~12 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[7]~12 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~12 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_mask[7]~q ),
	.datac(!\M_rot_pass3~q ),
	.datad(!\M_rot_sel_fill3~q ),
	.datae(!\M_rot[7]~12_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~12 .extended_lut = "off";
defparam \A_shift_rot_result~12 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~12 .shared_arith = "off";

dffeas \A_shift_rot_result[31] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~12_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_shift_rot_result[31]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[31] .is_wysiwyg = "true";
defparam \A_shift_rot_result[31] .power_up = "low";

dffeas \A_inst_result[31] (
	.clk(clk_clk),
	.d(\M_alu_result[31]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\A_inst_result[26]~1_combout ),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_inst_result[31]~q ),
	.prn(vcc));
defparam \A_inst_result[31] .is_wysiwyg = "true";
defparam \A_inst_result[31] .power_up = "low";

cyclonev_lcell_comb \Add11~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[15]~q ),
	.datae(gnd),
	.dataf(!\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[31]~q ),
	.datag(gnd),
	.cin(\Add11~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add11~17_sumout ),
	.cout(),
	.shareout());
defparam \Add11~17 .extended_lut = "off";
defparam \Add11~17 .lut_mask = 64'h0000FF00000000FF;
defparam \Add11~17 .shared_arith = "off";

dffeas \A_mul_s1[15] (
	.clk(clk_clk),
	.d(\Add11~17_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_mul_s1[15]~q ),
	.prn(vcc));
defparam \A_mul_s1[15] .is_wysiwyg = "true";
defparam \A_mul_s1[15] .power_up = "low";

dffeas \A_mul_cell_p3[15] (
	.clk(clk_clk),
	.d(\the_first_nios2_system_cpu_cpu_mult_cell|the_altmult_add_p3|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[15]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_mul_cell_p3[15]~q ),
	.prn(vcc));
defparam \A_mul_cell_p3[15] .is_wysiwyg = "true";
defparam \A_mul_cell_p3[15] .power_up = "low";

cyclonev_lcell_comb \Add12~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_mul_s1[15]~q ),
	.datae(gnd),
	.dataf(!\A_mul_cell_p3[15]~q ),
	.datag(gnd),
	.cin(\Add12~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add12~17_sumout ),
	.cout(),
	.shareout());
defparam \Add12~17 .extended_lut = "off";
defparam \Add12~17 .lut_mask = 64'h0000FF00000000FF;
defparam \Add12~17 .shared_arith = "off";

cyclonev_lcell_comb \A_wr_data_unfiltered[31]~14 (
	.dataa(!\A_slow_inst_result[31]~q ),
	.datab(!\A_shift_rot_result[31]~q ),
	.datac(!\A_inst_result[31]~q ),
	.datad(!\Add12~17_sumout ),
	.datae(!\A_wr_data_unfiltered[15]~0_combout ),
	.dataf(!\A_wr_data_unfiltered[15]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[31]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[31]~14 .extended_lut = "off";
defparam \A_wr_data_unfiltered[31]~14 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_wr_data_unfiltered[31]~14 .shared_arith = "off";

dffeas \W_wr_data[31] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[31]~14_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[31]~q ),
	.prn(vcc));
defparam \W_wr_data[31] .is_wysiwyg = "true";
defparam \W_wr_data[31] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[31]~7 (
	.dataa(!\M_alu_result[31]~q ),
	.datab(!\A_wr_data_unfiltered[31]~14_combout ),
	.datac(!\first_nios2_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[31] ),
	.datad(!\W_wr_data[31]~q ),
	.datae(!\E_src1[26]~0_combout ),
	.dataf(!\E_src1[26]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[31]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[31]~7 .extended_lut = "off";
defparam \D_src1_reg[31]~7 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[31]~7 .shared_arith = "off";

dffeas \E_src1[31] (
	.clk(clk_clk),
	.d(\D_src1_reg[31]~7_combout ),
	.asdata(\E_alu_result[31]~combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\Equal303~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(!\A_mem_stall~q ),
	.q(\E_src1[31]~q ),
	.prn(vcc));
defparam \E_src1[31] .is_wysiwyg = "true";
defparam \E_src1[31] .power_up = "low";

cyclonev_lcell_comb \Add9~73 (
	.dataa(!\E_ctrl_alu_signed_comparison~q ),
	.datab(!\E_ctrl_alu_subtract~q ),
	.datac(gnd),
	.datad(!\E_src2[31]~q ),
	.datae(gnd),
	.dataf(!\E_src1[31]~q ),
	.datag(gnd),
	.cin(\Add9~122 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~73_sumout ),
	.cout(\Add9~74 ),
	.shareout());
defparam \Add9~73 .extended_lut = "off";
defparam \Add9~73 .lut_mask = 64'h000055AA00009966;
defparam \Add9~73 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[31]~33 (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\D_src2_reg[0]~2_combout ),
	.datac(!\Add9~73_sumout ),
	.datad(!\E_alu_result~10_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[31]~33_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[31]~33 .extended_lut = "off";
defparam \D_src2_reg[31]~33 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \D_src2_reg[31]~33 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[31]~35 (
	.dataa(!\D_ctrl_b_is_dst~q ),
	.datab(!\A_regnum_b_cmp_D~q ),
	.datac(!\M_regnum_b_cmp_D~q ),
	.datad(!\W_wr_data[31]~q ),
	.datae(!\M_alu_result[31]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[31]~35_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[31]~35 .extended_lut = "off";
defparam \D_src2_reg[31]~35 .lut_mask = 64'hDEFFFFFFDEFFFFFF;
defparam \D_src2_reg[31]~35 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[31]~36 (
	.dataa(!\D_src2_reg[0]~9_combout ),
	.datab(!\D_src2_reg[27]~34_combout ),
	.datac(!\A_wr_data_unfiltered[31]~14_combout ),
	.datad(!\D_src2_reg[31]~35_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[31]~36_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[31]~36 .extended_lut = "off";
defparam \D_src2_reg[31]~36 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \D_src2_reg[31]~36 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[31]~9 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\D_ctrl_src2_choose_imm~q ),
	.datac(!\D_ctrl_shift_right_arith~0_combout ),
	.datad(!\D_iw[21]~q ),
	.datae(!\D_ctrl_unsigned_lo_imm16~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[31]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[31]~9 .extended_lut = "off";
defparam \D_src2[31]~9 .lut_mask = 64'hFFFFF7FFFFFFF7FF;
defparam \D_src2[31]~9 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[31]~10 (
	.dataa(!\D_src2_reg[0]~6_combout ),
	.datab(!\D_ctrl_src2_choose_imm~q ),
	.datac(!\D_src2_reg[31]~33_combout ),
	.datad(!\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[31] ),
	.datae(!\D_src2_reg[31]~36_combout ),
	.dataf(!\D_src2[31]~9_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[31]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[31]~10 .extended_lut = "off";
defparam \D_src2[31]~10 .lut_mask = 64'hDFFFFFFFFFFFFFFF;
defparam \D_src2[31]~10 .shared_arith = "off";

dffeas \E_src2[31] (
	.clk(clk_clk),
	.d(\D_src2[31]~10_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_src2[31]~q ),
	.prn(vcc));
defparam \E_src2[31] .is_wysiwyg = "true";
defparam \E_src2[31] .power_up = "low";

cyclonev_lcell_comb \Add9~61 (
	.dataa(gnd),
	.datab(!\E_ctrl_alu_subtract~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add9~74 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~61_sumout ),
	.cout(),
	.shareout());
defparam \Add9~61 .extended_lut = "off";
defparam \Add9~61 .lut_mask = 64'h0000000000003333;
defparam \Add9~61 .shared_arith = "off";

dffeas \E_bht_data[1] (
	.clk(clk_clk),
	.d(\D_bht_data[1]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_bht_data[1]~q ),
	.prn(vcc));
defparam \E_bht_data[1] .is_wysiwyg = "true";
defparam \E_bht_data[1] .power_up = "low";

dffeas E_ctrl_br_cond(
	.clk(clk_clk),
	.d(\E_ctrl_br_cond_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_ctrl_br_cond~q ),
	.prn(vcc));
defparam E_ctrl_br_cond.is_wysiwyg = "true";
defparam E_ctrl_br_cond.power_up = "low";

cyclonev_lcell_comb \E_br_mispredict~0 (
	.dataa(!\E_valid~combout ),
	.datab(!\E_ctrl_br_cond~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_br_mispredict~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_br_mispredict~0 .extended_lut = "off";
defparam \E_br_mispredict~0 .lut_mask = 64'h7777777777777777;
defparam \E_br_mispredict~0 .shared_arith = "off";

cyclonev_lcell_comb M_pipe_flush_nxt(
	.dataa(!\A_pipe_flush_nxt~0_combout ),
	.datab(!\Add9~61_sumout ),
	.datac(!\E_br_result~0_combout ),
	.datad(!\E_br_result~1_combout ),
	.datae(!\E_bht_data[1]~q ),
	.dataf(!\E_br_mispredict~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_pipe_flush_nxt~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam M_pipe_flush_nxt.extended_lut = "off";
defparam M_pipe_flush_nxt.lut_mask = 64'hFFFFFFFFBEEBEBBE;
defparam M_pipe_flush_nxt.shared_arith = "off";

dffeas M_pipe_flush(
	.clk(clk_clk),
	.d(\M_pipe_flush_nxt~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_pipe_flush~q ),
	.prn(vcc));
defparam M_pipe_flush.is_wysiwyg = "true";
defparam M_pipe_flush.power_up = "low";

cyclonev_lcell_comb \D_ctrl_shift_rot~1 (
	.dataa(!\D_iw[14]~q ),
	.datab(!\D_iw[13]~q ),
	.datac(!\D_iw[12]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_shift_rot~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_shift_rot~1 .extended_lut = "off";
defparam \D_ctrl_shift_rot~1 .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \D_ctrl_shift_rot~1 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_late_result~1 (
	.dataa(!\D_iw[16]~q ),
	.datab(!\D_iw[15]~q ),
	.datac(!\D_iw[14]~q ),
	.datad(!\D_iw[13]~q ),
	.datae(!\D_iw[12]~q ),
	.dataf(!\D_iw[11]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_late_result~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_late_result~1 .extended_lut = "off";
defparam \D_ctrl_late_result~1 .lut_mask = 64'hDDF5FFFFFFFFFFFF;
defparam \D_ctrl_late_result~1 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_late_result~0 (
	.dataa(!\Equal95~0_combout ),
	.datab(!\D_ctrl_ld~0_combout ),
	.datac(!\Equal95~7_combout ),
	.datad(!\D_ctrl_shift_rot~1_combout ),
	.datae(!\D_ctrl_late_result~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_late_result~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_late_result~0 .extended_lut = "off";
defparam \D_ctrl_late_result~0 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \D_ctrl_late_result~0 .shared_arith = "off";

dffeas E_ctrl_late_result(
	.clk(clk_clk),
	.d(\D_ctrl_late_result~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_ctrl_late_result~q ),
	.prn(vcc));
defparam E_ctrl_late_result.is_wysiwyg = "true";
defparam E_ctrl_late_result.power_up = "low";

cyclonev_lcell_comb \D_data_depend~0 (
	.dataa(!\D_ctrl_b_is_dst~q ),
	.datab(!\E_regnum_b_cmp_D~q ),
	.datac(!\E_ctrl_late_result~q ),
	.datad(!\D_ctrl_a_not_src~q ),
	.datae(!\E_regnum_a_cmp_D~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_data_depend~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_data_depend~0 .extended_lut = "off";
defparam \D_data_depend~0 .lut_mask = 64'hFFBFFFFFFFBFFFFF;
defparam \D_data_depend~0 .shared_arith = "off";

dffeas M_ctrl_late_result(
	.clk(clk_clk),
	.d(\E_ctrl_late_result~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_ctrl_late_result~q ),
	.prn(vcc));
defparam M_ctrl_late_result.is_wysiwyg = "true";
defparam M_ctrl_late_result.power_up = "low";

cyclonev_lcell_comb \D_data_depend~1 (
	.dataa(!\D_ctrl_b_is_dst~q ),
	.datab(!\M_regnum_b_cmp_D~q ),
	.datac(!\D_ctrl_a_not_src~q ),
	.datad(!\M_regnum_a_cmp_D~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_data_depend~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_data_depend~1 .extended_lut = "off";
defparam \D_data_depend~1 .lut_mask = 64'hFBFFFBFFFBFFFBFF;
defparam \D_data_depend~1 .shared_arith = "off";

cyclonev_lcell_comb D_valid(
	.dataa(!\M_pipe_flush~q ),
	.datab(!\D_issue~q ),
	.datac(!\D_data_depend~0_combout ),
	.datad(!\M_ctrl_late_result~q ),
	.datae(!\D_data_depend~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_valid~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam D_valid.extended_lut = "off";
defparam D_valid.lut_mask = 64'hFFFFFFF7FFFFFFF7;
defparam D_valid.shared_arith = "off";

dffeas E_valid_from_D(
	.clk(clk_clk),
	.d(\D_valid~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_valid_from_D~q ),
	.prn(vcc));
defparam E_valid_from_D.is_wysiwyg = "true";
defparam E_valid_from_D.power_up = "low";

cyclonev_lcell_comb E_valid(
	.dataa(!\E_valid_from_D~q ),
	.datab(!\M_pipe_flush~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_valid~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam E_valid.extended_lut = "off";
defparam E_valid.lut_mask = 64'h7777777777777777;
defparam E_valid.shared_arith = "off";

dffeas M_valid_from_E(
	.clk(clk_clk),
	.d(\E_valid~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_valid_from_E~q ),
	.prn(vcc));
defparam M_valid_from_E.is_wysiwyg = "true";
defparam M_valid_from_E.power_up = "low";

cyclonev_lcell_comb \M_exc_allowed~0 (
	.dataa(!\M_valid_from_E~q ),
	.datab(!\A_pipe_flush~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_exc_allowed~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_exc_allowed~0 .extended_lut = "off";
defparam \M_exc_allowed~0 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \M_exc_allowed~0 .shared_arith = "off";

dffeas A_exc_allowed(
	.clk(clk_clk),
	.d(\M_exc_allowed~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_exc_allowed~q ),
	.prn(vcc));
defparam A_exc_allowed.is_wysiwyg = "true";
defparam A_exc_allowed.power_up = "low";

cyclonev_lcell_comb \wait_for_one_post_bret_inst~1 (
	.dataa(!W_debug_mode1),
	.datab(!\the_first_nios2_system_cpu_cpu_nios2_oci|the_first_nios2_system_cpu_cpu_nios2_avalon_reg|oci_single_step_mode~q ),
	.datac(!\wait_for_one_post_bret_inst~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_for_one_post_bret_inst~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_for_one_post_bret_inst~1 .extended_lut = "off";
defparam \wait_for_one_post_bret_inst~1 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \wait_for_one_post_bret_inst~1 .shared_arith = "off";

dffeas wait_for_one_post_bret_inst(
	.clk(clk_clk),
	.d(\wait_for_one_post_bret_inst~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wait_for_one_post_bret_inst~q ),
	.prn(vcc));
defparam wait_for_one_post_bret_inst.is_wysiwyg = "true";
defparam wait_for_one_post_bret_inst.power_up = "low";

cyclonev_lcell_comb \wait_for_one_post_bret_inst~0 (
	.dataa(!\A_valid_from_M~q ),
	.datab(!\A_exc_any~q ),
	.datac(!\A_exc_allowed~q ),
	.datad(!\wait_for_one_post_bret_inst~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_for_one_post_bret_inst~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_for_one_post_bret_inst~0 .extended_lut = "off";
defparam \wait_for_one_post_bret_inst~0 .lut_mask = 64'hFEFFFEFFFEFFFEFF;
defparam \wait_for_one_post_bret_inst~0 .shared_arith = "off";

cyclonev_lcell_comb \hbreak_req~0 (
	.dataa(!W_debug_mode1),
	.datab(!\the_first_nios2_system_cpu_cpu_nios2_oci|the_first_nios2_system_cpu_cpu_nios2_avalon_reg|oci_single_step_mode~q ),
	.datac(!\wait_for_one_post_bret_inst~0_combout ),
	.datad(!\latched_oci_tb_hbreak_req~q ),
	.datae(!\the_first_nios2_system_cpu_cpu_nios2_oci|the_first_nios2_system_cpu_cpu_nios2_oci_debug|jtag_break~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\hbreak_req~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \hbreak_req~0 .extended_lut = "off";
defparam \hbreak_req~0 .lut_mask = 64'hFEFFFFFFFEFFFFFF;
defparam \hbreak_req~0 .shared_arith = "off";

cyclonev_lcell_comb M_exc_any(
	.dataa(!\M_norm_intr_req~q ),
	.datab(!\hbreak_req~0_combout ),
	.datac(!\M_exc_any~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_exc_any~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam M_exc_any.extended_lut = "off";
defparam M_exc_any.lut_mask = 64'hF7F7F7F7F7F7F7F7;
defparam M_exc_any.shared_arith = "off";

dffeas A_exc_any(
	.clk(clk_clk),
	.d(\M_exc_any~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_exc_any~q ),
	.prn(vcc));
defparam A_exc_any.is_wysiwyg = "true";
defparam A_exc_any.power_up = "low";

dffeas \M_iw[11] (
	.clk(clk_clk),
	.d(\E_iw[11]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_iw[11]~q ),
	.prn(vcc));
defparam \M_iw[11] .is_wysiwyg = "true";
defparam \M_iw[11] .power_up = "low";

dffeas \A_iw[11] (
	.clk(clk_clk),
	.d(\M_iw[11]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_iw[11]~q ),
	.prn(vcc));
defparam \A_iw[11] .is_wysiwyg = "true";
defparam \A_iw[11] .power_up = "low";

dffeas \M_iw[5] (
	.clk(clk_clk),
	.d(\E_iw[5]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_iw[5]~q ),
	.prn(vcc));
defparam \M_iw[5] .is_wysiwyg = "true";
defparam \M_iw[5] .power_up = "low";

dffeas \A_iw[5] (
	.clk(clk_clk),
	.d(\M_iw[5]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_iw[5]~q ),
	.prn(vcc));
defparam \A_iw[5] .is_wysiwyg = "true";
defparam \A_iw[5] .power_up = "low";

dffeas \M_iw[0] (
	.clk(clk_clk),
	.d(\E_iw[0]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_iw[0]~q ),
	.prn(vcc));
defparam \M_iw[0] .is_wysiwyg = "true";
defparam \M_iw[0] .power_up = "low";

dffeas \A_iw[0] (
	.clk(clk_clk),
	.d(\M_iw[0]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_iw[0]~q ),
	.prn(vcc));
defparam \A_iw[0] .is_wysiwyg = "true";
defparam \A_iw[0] .power_up = "low";

dffeas \M_iw[16] (
	.clk(clk_clk),
	.d(\E_iw[16]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_iw[16]~q ),
	.prn(vcc));
defparam \M_iw[16] .is_wysiwyg = "true";
defparam \M_iw[16] .power_up = "low";

dffeas \A_iw[16] (
	.clk(clk_clk),
	.d(\M_iw[16]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_iw[16]~q ),
	.prn(vcc));
defparam \A_iw[16] .is_wysiwyg = "true";
defparam \A_iw[16] .power_up = "low";

dffeas \M_iw[15] (
	.clk(clk_clk),
	.d(\E_iw[15]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_iw[15]~q ),
	.prn(vcc));
defparam \M_iw[15] .is_wysiwyg = "true";
defparam \M_iw[15] .power_up = "low";

dffeas \A_iw[15] (
	.clk(clk_clk),
	.d(\M_iw[15]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_iw[15]~q ),
	.prn(vcc));
defparam \A_iw[15] .is_wysiwyg = "true";
defparam \A_iw[15] .power_up = "low";

dffeas \M_iw[13] (
	.clk(clk_clk),
	.d(\E_iw[13]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_iw[13]~q ),
	.prn(vcc));
defparam \M_iw[13] .is_wysiwyg = "true";
defparam \M_iw[13] .power_up = "low";

dffeas \A_iw[13] (
	.clk(clk_clk),
	.d(\M_iw[13]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_iw[13]~q ),
	.prn(vcc));
defparam \A_iw[13] .is_wysiwyg = "true";
defparam \A_iw[13] .power_up = "low";

dffeas \M_iw[12] (
	.clk(clk_clk),
	.d(\E_iw[12]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_iw[12]~q ),
	.prn(vcc));
defparam \M_iw[12] .is_wysiwyg = "true";
defparam \M_iw[12] .power_up = "low";

dffeas \A_iw[12] (
	.clk(clk_clk),
	.d(\M_iw[12]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_iw[12]~q ),
	.prn(vcc));
defparam \A_iw[12] .is_wysiwyg = "true";
defparam \A_iw[12] .power_up = "low";

cyclonev_lcell_comb \A_op_eret~0 (
	.dataa(!\A_iw[16]~q ),
	.datab(!\A_iw[15]~q ),
	.datac(!\A_iw[13]~q ),
	.datad(!\A_iw[12]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_op_eret~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_op_eret~0 .extended_lut = "off";
defparam \A_op_eret~0 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \A_op_eret~0 .shared_arith = "off";

dffeas \M_iw[4] (
	.clk(clk_clk),
	.d(\E_iw[4]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_iw[4]~q ),
	.prn(vcc));
defparam \M_iw[4] .is_wysiwyg = "true";
defparam \M_iw[4] .power_up = "low";

dffeas \A_iw[4] (
	.clk(clk_clk),
	.d(\M_iw[4]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_iw[4]~q ),
	.prn(vcc));
defparam \A_iw[4] .is_wysiwyg = "true";
defparam \A_iw[4] .power_up = "low";

dffeas \M_iw[3] (
	.clk(clk_clk),
	.d(\E_iw[3]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_iw[3]~q ),
	.prn(vcc));
defparam \M_iw[3] .is_wysiwyg = "true";
defparam \M_iw[3] .power_up = "low";

dffeas \A_iw[3] (
	.clk(clk_clk),
	.d(\M_iw[3]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_iw[3]~q ),
	.prn(vcc));
defparam \A_iw[3] .is_wysiwyg = "true";
defparam \A_iw[3] .power_up = "low";

dffeas \M_iw[2] (
	.clk(clk_clk),
	.d(\E_iw[2]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_iw[2]~q ),
	.prn(vcc));
defparam \M_iw[2] .is_wysiwyg = "true";
defparam \M_iw[2] .power_up = "low";

dffeas \A_iw[2] (
	.clk(clk_clk),
	.d(\M_iw[2]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_iw[2]~q ),
	.prn(vcc));
defparam \A_iw[2] .is_wysiwyg = "true";
defparam \A_iw[2] .power_up = "low";

dffeas \M_iw[1] (
	.clk(clk_clk),
	.d(\E_iw[1]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_iw[1]~q ),
	.prn(vcc));
defparam \M_iw[1] .is_wysiwyg = "true";
defparam \M_iw[1] .power_up = "low";

dffeas \A_iw[1] (
	.clk(clk_clk),
	.d(\M_iw[1]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_iw[1]~q ),
	.prn(vcc));
defparam \A_iw[1] .is_wysiwyg = "true";
defparam \A_iw[1] .power_up = "low";

cyclonev_lcell_comb \A_op_eret~1 (
	.dataa(!\A_iw[4]~q ),
	.datab(!\A_iw[3]~q ),
	.datac(!\A_iw[2]~q ),
	.datad(!\A_iw[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_op_eret~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_op_eret~1 .extended_lut = "off";
defparam \A_op_eret~1 .lut_mask = 64'hF7FFF7FFF7FFF7FF;
defparam \A_op_eret~1 .shared_arith = "off";

cyclonev_lcell_comb \A_op_eret~2 (
	.dataa(!\A_iw[11]~q ),
	.datab(!\A_iw[5]~q ),
	.datac(!\A_iw[0]~q ),
	.datad(!\A_op_eret~0_combout ),
	.datae(!\A_op_eret~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_op_eret~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_op_eret~2 .extended_lut = "off";
defparam \A_op_eret~2 .lut_mask = 64'hF7FFFFFFF7FFFFFF;
defparam \A_op_eret~2 .shared_arith = "off";

cyclonev_lcell_comb \W_status_reg_pie_nxt~0 (
	.dataa(gnd),
	.datab(!\A_op_eret~2_combout ),
	.datac(!\A_iw[7]~q ),
	.datad(!\A_iw[6]~q ),
	.datae(!\A_wrctl_status~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_status_reg_pie_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_status_reg_pie_nxt~0 .extended_lut = "off";
defparam \W_status_reg_pie_nxt~0 .lut_mask = 64'hFFFFCFFFFFFFCFFF;
defparam \W_status_reg_pie_nxt~0 .shared_arith = "off";

dffeas \M_iw[14] (
	.clk(clk_clk),
	.d(\E_iw[14]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_iw[14]~q ),
	.prn(vcc));
defparam \M_iw[14] .is_wysiwyg = "true";
defparam \M_iw[14] .power_up = "low";

dffeas \A_iw[14] (
	.clk(clk_clk),
	.d(\M_iw[14]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_iw[14]~q ),
	.prn(vcc));
defparam \A_iw[14] .is_wysiwyg = "true";
defparam \A_iw[14] .power_up = "low";

cyclonev_lcell_comb \W_status_reg_pie_nxt~1 (
	.dataa(!\A_inst_result[0]~q ),
	.datab(!\A_iw[7]~q ),
	.datac(!\A_iw[6]~q ),
	.datad(!\A_wrctl_status~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_status_reg_pie_nxt~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_status_reg_pie_nxt~1 .extended_lut = "off";
defparam \W_status_reg_pie_nxt~1 .lut_mask = 64'hFDFFFDFFFDFFFDFF;
defparam \W_status_reg_pie_nxt~1 .shared_arith = "off";

cyclonev_lcell_comb \W_status_reg_pie_nxt~2 (
	.dataa(!\A_iw[14]~q ),
	.datab(!\A_op_eret~2_combout ),
	.datac(!\W_estatus_reg_pie~q ),
	.datad(!\W_bstatus_reg_pie~q ),
	.datae(!\W_status_reg_pie_nxt~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_status_reg_pie_nxt~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_status_reg_pie_nxt~2 .extended_lut = "off";
defparam \W_status_reg_pie_nxt~2 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \W_status_reg_pie_nxt~2 .shared_arith = "off";

cyclonev_lcell_comb \W_status_reg_pie_nxt~3 (
	.dataa(!\A_valid_from_M~q ),
	.datab(!\A_exc_any~q ),
	.datac(!\A_exc_allowed~q ),
	.datad(!\W_status_reg_pie~q ),
	.datae(!\W_status_reg_pie_nxt~0_combout ),
	.dataf(!\W_status_reg_pie_nxt~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_status_reg_pie_nxt~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_status_reg_pie_nxt~3 .extended_lut = "off";
defparam \W_status_reg_pie_nxt~3 .lut_mask = 64'hD8FFFFFFFFFFFFFF;
defparam \W_status_reg_pie_nxt~3 .shared_arith = "off";

dffeas W_status_reg_pie(
	.clk(clk_clk),
	.d(\W_status_reg_pie_nxt~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_status_reg_pie~q ),
	.prn(vcc));
defparam W_status_reg_pie.is_wysiwyg = "true";
defparam W_status_reg_pie.power_up = "low";

cyclonev_lcell_comb \norm_intr_req~0 (
	.dataa(!\W_status_reg_pie~q ),
	.datab(!\W_ipending_reg_irq1~q ),
	.datac(!\W_ipending_reg_irq16~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\norm_intr_req~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \norm_intr_req~0 .extended_lut = "off";
defparam \norm_intr_req~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \norm_intr_req~0 .shared_arith = "off";

dffeas M_norm_intr_req(
	.clk(clk_clk),
	.d(\norm_intr_req~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_norm_intr_req~q ),
	.prn(vcc));
defparam M_norm_intr_req.is_wysiwyg = "true";
defparam M_norm_intr_req.power_up = "low";

cyclonev_lcell_comb \M_valid~0 (
	.dataa(!\M_norm_intr_req~q ),
	.datab(!\hbreak_req~0_combout ),
	.datac(!\M_exc_allowed~0_combout ),
	.datad(!\M_exc_any~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_valid~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_valid~0 .extended_lut = "off";
defparam \M_valid~0 .lut_mask = 64'hEFFFEFFFEFFFEFFF;
defparam \M_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \M_data_master_start_stall~0 (
	.dataa(!\A_mem_stall~q ),
	.datab(!\M_sel_data_master~q ),
	.datac(!\M_valid~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_data_master_start_stall~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_data_master_start_stall~0 .extended_lut = "off";
defparam \M_data_master_start_stall~0 .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \M_data_master_start_stall~0 .shared_arith = "off";

cyclonev_lcell_comb \E_ctrl_ld_st~0 (
	.dataa(!\E_iw[1]~q ),
	.datab(!\E_iw[2]~q ),
	.datac(!\E_iw[4]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_ctrl_ld_st~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_ctrl_ld_st~0 .extended_lut = "off";
defparam \E_ctrl_ld_st~0 .lut_mask = 64'hF7F7F7F7F7F7F7F7;
defparam \E_ctrl_ld_st~0 .shared_arith = "off";

dffeas M_ctrl_ld_st(
	.clk(clk_clk),
	.d(\E_ctrl_ld_st~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(!\E_iw[0]~q ),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_ctrl_ld_st~q ),
	.prn(vcc));
defparam M_ctrl_ld_st.is_wysiwyg = "true";
defparam M_ctrl_ld_st.power_up = "low";

cyclonev_lcell_comb \E_ctrl_st~0 (
	.dataa(!\E_iw[1]~q ),
	.datab(!\E_iw[2]~q ),
	.datac(!\E_iw[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_ctrl_st~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_ctrl_st~0 .extended_lut = "off";
defparam \E_ctrl_st~0 .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \E_ctrl_st~0 .shared_arith = "off";

dffeas M_ctrl_st(
	.clk(clk_clk),
	.d(\E_ctrl_st~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_ctrl_st~q ),
	.prn(vcc));
defparam M_ctrl_st.is_wysiwyg = "true";
defparam M_ctrl_st.power_up = "low";

dffeas A_ctrl_st(
	.clk(clk_clk),
	.d(\M_ctrl_st~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_ctrl_st~q ),
	.prn(vcc));
defparam A_ctrl_st.is_wysiwyg = "true";
defparam A_ctrl_st.power_up = "low";

cyclonev_lcell_comb M_data_master_start_stall(
	.dataa(!\M_data_master_start_stall~0_combout ),
	.datab(!\M_ctrl_ld_st~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_data_master_start_stall~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam M_data_master_start_stall.extended_lut = "off";
defparam M_data_master_start_stall.lut_mask = 64'h7777777777777777;
defparam M_data_master_start_stall.shared_arith = "off";

dffeas A_data_master_started_stall(
	.clk(clk_clk),
	.d(\M_data_master_start_stall~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_data_master_started_stall~q ),
	.prn(vcc));
defparam A_data_master_started_stall.is_wysiwyg = "true";
defparam A_data_master_started_stall.power_up = "low";

cyclonev_lcell_comb \av_ld_data_transfer~0 (
	.dataa(!d_read1),
	.datab(!read_latency_shift_reg_0),
	.datac(!WideOr1),
	.datad(!WideOr11),
	.datae(!WideOr12),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_data_transfer~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_data_transfer~0 .extended_lut = "off";
defparam \av_ld_data_transfer~0 .lut_mask = 64'hFFFFFFF7FFFFFFF7;
defparam \av_ld_data_transfer~0 .shared_arith = "off";

dffeas av_ld_aligning_data(
	.clk(clk_clk),
	.d(\av_ld_data_transfer~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\av_ld_aligning_data~q ),
	.prn(vcc));
defparam av_ld_aligning_data.is_wysiwyg = "true";
defparam av_ld_aligning_data.power_up = "low";

cyclonev_lcell_comb \A_mem_stall_nxt~0 (
	.dataa(!\A_data_master_started_stall~q ),
	.datab(!\A_ctrl_st~q ),
	.datac(!\av_ld_aligning_data~q ),
	.datad(!\A_ctrl_ld32~q ),
	.datae(!\av_ld_data_transfer~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_mem_stall_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_mem_stall_nxt~0 .extended_lut = "off";
defparam \A_mem_stall_nxt~0 .lut_mask = 64'h5F3FFFFF5F3FFFFF;
defparam \A_mem_stall_nxt~0 .shared_arith = "off";

cyclonev_lcell_comb \A_mem_stall_nxt~1 (
	.dataa(!\A_mem_stall~q ),
	.datab(!\M_data_master_start_stall~0_combout ),
	.datac(!av_waitrequest),
	.datad(!\M_ctrl_ld_st~q ),
	.datae(!\A_ctrl_st~q ),
	.dataf(!\A_mem_stall_nxt~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_mem_stall_nxt~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_mem_stall_nxt~1 .extended_lut = "off";
defparam \A_mem_stall_nxt~1 .lut_mask = 64'hF7FFFFFFB3FFFFFF;
defparam \A_mem_stall_nxt~1 .shared_arith = "off";

dffeas A_mem_stall(
	.clk(clk_clk),
	.d(\A_mem_stall_nxt~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mem_stall~q ),
	.prn(vcc));
defparam A_mem_stall.is_wysiwyg = "true";
defparam A_mem_stall.power_up = "low";

cyclonev_lcell_comb \F_stall~0 (
	.dataa(!\A_mem_stall~q ),
	.datab(!\M_pipe_flush~q ),
	.datac(!\D_issue~q ),
	.datad(!\D_data_depend~0_combout ),
	.datae(!\M_ctrl_late_result~q ),
	.dataf(!\D_data_depend~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_stall~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_stall~0 .extended_lut = "off";
defparam \F_stall~0 .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \F_stall~0 .shared_arith = "off";

dffeas \D_iw[5] (
	.clk(clk_clk),
	.d(\first_nios2_system_cpu_cpu_ic_data|the_altsyncram|auto_generated|q_b[5] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_iw[5]~q ),
	.prn(vcc));
defparam \D_iw[5] .is_wysiwyg = "true";
defparam \D_iw[5] .power_up = "low";

cyclonev_lcell_comb \D_ctrl_cmp~0 (
	.dataa(!\D_iw[5]~q ),
	.datab(!\D_iw[4]~q ),
	.datac(!\D_iw[3]~q ),
	.datad(!\D_iw[2]~q ),
	.datae(!\D_iw[1]~q ),
	.dataf(!\D_iw[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_cmp~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_cmp~0 .extended_lut = "off";
defparam \D_ctrl_cmp~0 .lut_mask = 64'hFFFFFFFFFFFFFF96;
defparam \D_ctrl_cmp~0 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_cmp~1 (
	.dataa(!\D_iw[5]~q ),
	.datab(!\D_iw[4]~q ),
	.datac(!\D_iw[3]~q ),
	.datad(!\D_iw[2]~q ),
	.datae(!\D_iw[1]~q ),
	.dataf(!\D_iw[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_cmp~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_cmp~1 .extended_lut = "off";
defparam \D_ctrl_cmp~1 .lut_mask = 64'hFFFFFFFFFF69FF96;
defparam \D_ctrl_cmp~1 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_cmp~3 (
	.dataa(!\D_iw[13]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[11]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_cmp~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_cmp~3 .extended_lut = "off";
defparam \D_ctrl_cmp~3 .lut_mask = 64'hFEFEFEFEFEFEFEFE;
defparam \D_ctrl_cmp~3 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_cmp~2 (
	.dataa(!\D_ctrl_cmp~0_combout ),
	.datab(!\D_ctrl_cmp~1_combout ),
	.datac(gnd),
	.datad(!\D_ctrl_cmp~3_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_cmp~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_cmp~2 .extended_lut = "off";
defparam \D_ctrl_cmp~2 .lut_mask = 64'h5533553355335533;
defparam \D_ctrl_cmp~2 .shared_arith = "off";

dffeas E_ctrl_cmp(
	.clk(clk_clk),
	.d(\D_ctrl_cmp~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_ctrl_cmp~q ),
	.prn(vcc));
defparam E_ctrl_cmp.is_wysiwyg = "true";
defparam E_ctrl_cmp.power_up = "low";

cyclonev_lcell_comb \D_src2_reg[0]~3 (
	.dataa(!\E_ctrl_cmp~q ),
	.datab(!\Add9~61_sumout ),
	.datac(!\E_br_result~0_combout ),
	.datad(!\E_br_result~1_combout ),
	.datae(!\D_src2_reg[0]~2_combout ),
	.dataf(!\E_alu_result[0]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[0]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[0]~3 .extended_lut = "off";
defparam \D_src2_reg[0]~3 .lut_mask = 64'h47FFFFFFFFFFFFFF;
defparam \D_src2_reg[0]~3 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[0]~11 (
	.dataa(!\D_src2_reg[0]~3_combout ),
	.datab(!\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[0] ),
	.datac(!\D_src2_reg[0]~6_combout ),
	.datad(!\D_src2_reg[0]~10_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[0]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[0]~11 .extended_lut = "off";
defparam \D_src2_reg[0]~11 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \D_src2_reg[0]~11 .shared_arith = "off";

dffeas \E_src2_reg[0] (
	.clk(clk_clk),
	.d(\D_src2_reg[0]~11_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_src2_reg[0]~q ),
	.prn(vcc));
defparam \E_src2_reg[0] .is_wysiwyg = "true";
defparam \E_src2_reg[0] .power_up = "low";

dffeas \M_st_data[0] (
	.clk(clk_clk),
	.d(\E_src2_reg[0]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_st_data[0]~q ),
	.prn(vcc));
defparam \M_st_data[0] .is_wysiwyg = "true";
defparam \M_st_data[0] .power_up = "low";

dffeas \M_mem_baddr[4] (
	.clk(clk_clk),
	.d(\Add9~1_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_mem_baddr[4]~q ),
	.prn(vcc));
defparam \M_mem_baddr[4] .is_wysiwyg = "true";
defparam \M_mem_baddr[4] .power_up = "low";

dffeas \M_mem_baddr[5] (
	.clk(clk_clk),
	.d(\Add9~5_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_mem_baddr[5]~q ),
	.prn(vcc));
defparam \M_mem_baddr[5] .is_wysiwyg = "true";
defparam \M_mem_baddr[5] .power_up = "low";

dffeas \M_mem_baddr[8] (
	.clk(clk_clk),
	.d(\Add9~9_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_mem_baddr[8]~q ),
	.prn(vcc));
defparam \M_mem_baddr[8] .is_wysiwyg = "true";
defparam \M_mem_baddr[8] .power_up = "low";

dffeas \M_mem_baddr[16] (
	.clk(clk_clk),
	.d(\Add9~13_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_mem_baddr[16]~q ),
	.prn(vcc));
defparam \M_mem_baddr[16] .is_wysiwyg = "true";
defparam \M_mem_baddr[16] .power_up = "low";

dffeas \M_mem_baddr[15] (
	.clk(clk_clk),
	.d(\Add9~17_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_mem_baddr[15]~q ),
	.prn(vcc));
defparam \M_mem_baddr[15] .is_wysiwyg = "true";
defparam \M_mem_baddr[15] .power_up = "low";

dffeas \M_mem_baddr[14] (
	.clk(clk_clk),
	.d(\Add9~21_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_mem_baddr[14]~q ),
	.prn(vcc));
defparam \M_mem_baddr[14] .is_wysiwyg = "true";
defparam \M_mem_baddr[14] .power_up = "low";

dffeas \M_mem_baddr[13] (
	.clk(clk_clk),
	.d(\Add9~25_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_mem_baddr[13]~q ),
	.prn(vcc));
defparam \M_mem_baddr[13] .is_wysiwyg = "true";
defparam \M_mem_baddr[13] .power_up = "low";

dffeas \M_mem_baddr[12] (
	.clk(clk_clk),
	.d(\Add9~29_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_mem_baddr[12]~q ),
	.prn(vcc));
defparam \M_mem_baddr[12] .is_wysiwyg = "true";
defparam \M_mem_baddr[12] .power_up = "low";

dffeas \M_mem_baddr[11] (
	.clk(clk_clk),
	.d(\Add9~33_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_mem_baddr[11]~q ),
	.prn(vcc));
defparam \M_mem_baddr[11] .is_wysiwyg = "true";
defparam \M_mem_baddr[11] .power_up = "low";

dffeas \M_mem_baddr[10] (
	.clk(clk_clk),
	.d(\Add9~37_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_mem_baddr[10]~q ),
	.prn(vcc));
defparam \M_mem_baddr[10] .is_wysiwyg = "true";
defparam \M_mem_baddr[10] .power_up = "low";

dffeas \M_mem_baddr[9] (
	.clk(clk_clk),
	.d(\Add9~41_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_mem_baddr[9]~q ),
	.prn(vcc));
defparam \M_mem_baddr[9] .is_wysiwyg = "true";
defparam \M_mem_baddr[9] .power_up = "low";

dffeas \M_mem_baddr[7] (
	.clk(clk_clk),
	.d(\Add9~45_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_mem_baddr[7]~q ),
	.prn(vcc));
defparam \M_mem_baddr[7] .is_wysiwyg = "true";
defparam \M_mem_baddr[7] .power_up = "low";

dffeas \M_mem_baddr[6] (
	.clk(clk_clk),
	.d(\Add9~49_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_mem_baddr[6]~q ),
	.prn(vcc));
defparam \M_mem_baddr[6] .is_wysiwyg = "true";
defparam \M_mem_baddr[6] .power_up = "low";

cyclonev_lcell_comb d_write_nxt(
	.dataa(!d_write1),
	.datab(!\M_ctrl_st~q ),
	.datac(!\M_data_master_start_stall~0_combout ),
	.datad(!av_waitrequest),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_write_nxt~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam d_write_nxt.extended_lut = "off";
defparam d_write_nxt.lut_mask = 64'hFF7FFF7FFF7FFF7F;
defparam d_write_nxt.shared_arith = "off";

dffeas \M_mem_baddr[3] (
	.clk(clk_clk),
	.d(\Add9~53_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_mem_baddr[3]~q ),
	.prn(vcc));
defparam \M_mem_baddr[3] .is_wysiwyg = "true";
defparam \M_mem_baddr[3] .power_up = "low";

dffeas \M_mem_baddr[2] (
	.clk(clk_clk),
	.d(\Add9~57_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_mem_baddr[2]~q ),
	.prn(vcc));
defparam \M_mem_baddr[2] .is_wysiwyg = "true";
defparam \M_mem_baddr[2] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[1]~13 (
	.dataa(!\D_src2_reg[0]~4_combout ),
	.datab(!\D_src2_reg[0]~5_combout ),
	.datac(!\D_src2_reg[1]~12_combout ),
	.datad(!\E_alu_result[1]~combout ),
	.datae(!\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[1] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[1]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[1]~13 .extended_lut = "off";
defparam \D_src2_reg[1]~13 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \D_src2_reg[1]~13 .shared_arith = "off";

dffeas \E_src2_reg[1] (
	.clk(clk_clk),
	.d(\D_src2_reg[1]~13_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_src2_reg[1]~q ),
	.prn(vcc));
defparam \E_src2_reg[1] .is_wysiwyg = "true";
defparam \E_src2_reg[1] .power_up = "low";

dffeas \M_st_data[1] (
	.clk(clk_clk),
	.d(\E_src2_reg[1]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_st_data[1]~q ),
	.prn(vcc));
defparam \M_st_data[1] .is_wysiwyg = "true";
defparam \M_st_data[1] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[2]~15 (
	.dataa(!\D_src2_reg[0]~4_combout ),
	.datab(!\D_src2_reg[0]~5_combout ),
	.datac(!\D_src2_reg[2]~14_combout ),
	.datad(!\E_alu_result[2]~combout ),
	.datae(!\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[2] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[2]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[2]~15 .extended_lut = "off";
defparam \D_src2_reg[2]~15 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \D_src2_reg[2]~15 .shared_arith = "off";

dffeas \E_src2_reg[2] (
	.clk(clk_clk),
	.d(\D_src2_reg[2]~15_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_src2_reg[2]~q ),
	.prn(vcc));
defparam \E_src2_reg[2] .is_wysiwyg = "true";
defparam \E_src2_reg[2] .power_up = "low";

dffeas \M_st_data[2] (
	.clk(clk_clk),
	.d(\E_src2_reg[2]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_st_data[2]~q ),
	.prn(vcc));
defparam \M_st_data[2] .is_wysiwyg = "true";
defparam \M_st_data[2] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[3]~17 (
	.dataa(!\D_src2_reg[0]~4_combout ),
	.datab(!\D_src2_reg[0]~5_combout ),
	.datac(!\D_src2_reg[3]~16_combout ),
	.datad(!\E_alu_result[3]~combout ),
	.datae(!\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[3] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[3]~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[3]~17 .extended_lut = "off";
defparam \D_src2_reg[3]~17 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \D_src2_reg[3]~17 .shared_arith = "off";

dffeas \E_src2_reg[3] (
	.clk(clk_clk),
	.d(\D_src2_reg[3]~17_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_src2_reg[3]~q ),
	.prn(vcc));
defparam \E_src2_reg[3] .is_wysiwyg = "true";
defparam \E_src2_reg[3] .power_up = "low";

dffeas \M_st_data[3] (
	.clk(clk_clk),
	.d(\E_src2_reg[3]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_st_data[3]~q ),
	.prn(vcc));
defparam \M_st_data[3] .is_wysiwyg = "true";
defparam \M_st_data[3] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[4]~19 (
	.dataa(!\D_src2_reg[0]~4_combout ),
	.datab(!\D_src2_reg[0]~5_combout ),
	.datac(!\D_src2_reg[4]~18_combout ),
	.datad(!\E_alu_result[4]~combout ),
	.datae(!\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[4] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[4]~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[4]~19 .extended_lut = "off";
defparam \D_src2_reg[4]~19 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \D_src2_reg[4]~19 .shared_arith = "off";

dffeas \E_src2_reg[4] (
	.clk(clk_clk),
	.d(\D_src2_reg[4]~19_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_src2_reg[4]~q ),
	.prn(vcc));
defparam \E_src2_reg[4] .is_wysiwyg = "true";
defparam \E_src2_reg[4] .power_up = "low";

dffeas \M_st_data[4] (
	.clk(clk_clk),
	.d(\E_src2_reg[4]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_st_data[4]~q ),
	.prn(vcc));
defparam \M_st_data[4] .is_wysiwyg = "true";
defparam \M_st_data[4] .power_up = "low";

dffeas \E_src2_reg[5] (
	.clk(clk_clk),
	.d(\D_src2_reg[5]~21_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_src2_reg[5]~q ),
	.prn(vcc));
defparam \E_src2_reg[5] .is_wysiwyg = "true";
defparam \E_src2_reg[5] .power_up = "low";

dffeas \M_st_data[5] (
	.clk(clk_clk),
	.d(\E_src2_reg[5]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_st_data[5]~q ),
	.prn(vcc));
defparam \M_st_data[5] .is_wysiwyg = "true";
defparam \M_st_data[5] .power_up = "low";

dffeas \E_src2_reg[6] (
	.clk(clk_clk),
	.d(\D_src2_reg[6]~23_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_src2_reg[6]~q ),
	.prn(vcc));
defparam \E_src2_reg[6] .is_wysiwyg = "true";
defparam \E_src2_reg[6] .power_up = "low";

dffeas \M_st_data[6] (
	.clk(clk_clk),
	.d(\E_src2_reg[6]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_st_data[6]~q ),
	.prn(vcc));
defparam \M_st_data[6] .is_wysiwyg = "true";
defparam \M_st_data[6] .power_up = "low";

dffeas \E_src2_reg[7] (
	.clk(clk_clk),
	.d(\D_src2_reg[7]~25_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_src2_reg[7]~q ),
	.prn(vcc));
defparam \E_src2_reg[7] .is_wysiwyg = "true";
defparam \E_src2_reg[7] .power_up = "low";

dffeas \M_st_data[7] (
	.clk(clk_clk),
	.d(\E_src2_reg[7]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_st_data[7]~q ),
	.prn(vcc));
defparam \M_st_data[7] .is_wysiwyg = "true";
defparam \M_st_data[7] .power_up = "low";

cyclonev_lcell_comb d_read_nxt(
	.dataa(!d_read1),
	.datab(!\M_data_master_start_stall~0_combout ),
	.datac(!WideOr13),
	.datad(!\M_ctrl_ld~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_read_nxt~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam d_read_nxt.extended_lut = "off";
defparam d_read_nxt.lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam d_read_nxt.shared_arith = "off";

cyclonev_lcell_comb \W_debug_mode_nxt~0 (
	.dataa(!W_debug_mode1),
	.datab(!\A_valid_from_M~q ),
	.datac(!\A_exc_allowed~q ),
	.datad(!\A_exc_break~q ),
	.datae(!\A_iw[14]~q ),
	.dataf(!\A_op_eret~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_debug_mode_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_debug_mode_nxt~0 .extended_lut = "off";
defparam \W_debug_mode_nxt~0 .lut_mask = 64'hFFFFFFFFFFFFDFFF;
defparam \W_debug_mode_nxt~0 .shared_arith = "off";

cyclonev_lcell_comb \F_ic_fill_same_tag_line~0 (
	.dataa(!ic_fill_line_4),
	.datab(!ic_fill_line_3),
	.datac(!\F_pc[6]~q ),
	.datad(!\F_pc[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_fill_same_tag_line~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_fill_same_tag_line~0 .extended_lut = "off";
defparam \F_ic_fill_same_tag_line~0 .lut_mask = 64'h6996699669966996;
defparam \F_ic_fill_same_tag_line~0 .shared_arith = "off";

cyclonev_lcell_comb \F_ic_fill_same_tag_line~1 (
	.dataa(!ic_fill_line_1),
	.datab(!ic_fill_line_0),
	.datac(!\F_pc[3]~q ),
	.datad(!\F_pc[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_fill_same_tag_line~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_fill_same_tag_line~1 .extended_lut = "off";
defparam \F_ic_fill_same_tag_line~1 .lut_mask = 64'h6996699669966996;
defparam \F_ic_fill_same_tag_line~1 .shared_arith = "off";

cyclonev_lcell_comb \F_ic_fill_same_tag_line~2 (
	.dataa(!ic_fill_tag_1),
	.datab(!ic_fill_tag_0),
	.datac(!\F_pc[9]~q ),
	.datad(!\F_pc[10]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_fill_same_tag_line~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_fill_same_tag_line~2 .extended_lut = "off";
defparam \F_ic_fill_same_tag_line~2 .lut_mask = 64'h6996699669966996;
defparam \F_ic_fill_same_tag_line~2 .shared_arith = "off";

cyclonev_lcell_comb \F_ic_fill_same_tag_line~3 (
	.dataa(!ic_fill_tag_4),
	.datab(!ic_fill_tag_3),
	.datac(!\F_pc[12]~q ),
	.datad(!\F_pc[13]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_fill_same_tag_line~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_fill_same_tag_line~3 .extended_lut = "off";
defparam \F_ic_fill_same_tag_line~3 .lut_mask = 64'h6996699669966996;
defparam \F_ic_fill_same_tag_line~3 .shared_arith = "off";

cyclonev_lcell_comb \F_ic_fill_same_tag_line~4 (
	.dataa(!ic_fill_tag_5),
	.datab(!ic_fill_tag_2),
	.datac(!\F_pc[11]~q ),
	.datad(!\F_pc[14]~q ),
	.datae(!\F_ic_fill_same_tag_line~2_combout ),
	.dataf(!\F_ic_fill_same_tag_line~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_fill_same_tag_line~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_fill_same_tag_line~4 .extended_lut = "off";
defparam \F_ic_fill_same_tag_line~4 .lut_mask = 64'h6996FFFFFFFFFFFF;
defparam \F_ic_fill_same_tag_line~4 .shared_arith = "off";

cyclonev_lcell_comb \F_ic_fill_same_tag_line~5 (
	.dataa(!ic_fill_line_2),
	.datab(!\F_pc[5]~q ),
	.datac(!\F_ic_fill_same_tag_line~1_combout ),
	.datad(!\F_ic_fill_same_tag_line~4_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_fill_same_tag_line~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_fill_same_tag_line~5 .extended_lut = "off";
defparam \F_ic_fill_same_tag_line~5 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \F_ic_fill_same_tag_line~5 .shared_arith = "off";

cyclonev_lcell_comb F_ic_fill_same_tag_line(
	.dataa(!ic_fill_line_5),
	.datab(!\F_pc[8]~q ),
	.datac(!\F_ic_fill_same_tag_line~0_combout ),
	.datad(!\F_ic_fill_same_tag_line~5_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_fill_same_tag_line~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam F_ic_fill_same_tag_line.extended_lut = "off";
defparam F_ic_fill_same_tag_line.lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam F_ic_fill_same_tag_line.shared_arith = "off";

dffeas D_ic_fill_same_tag_line(
	.clk(clk_clk),
	.d(\F_ic_fill_same_tag_line~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~0_combout ),
	.q(\D_ic_fill_same_tag_line~q ),
	.prn(vcc));
defparam D_ic_fill_same_tag_line.is_wysiwyg = "true";
defparam D_ic_fill_same_tag_line.power_up = "low";

cyclonev_lcell_comb \E_ctrl_invalidate_i~0 (
	.dataa(!\E_iw[15]~q ),
	.datab(!\E_iw[12]~q ),
	.datac(!\E_iw[11]~q ),
	.datad(!\E_iw[16]~q ),
	.datae(!\E_iw[13]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_ctrl_invalidate_i~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_ctrl_invalidate_i~0 .extended_lut = "off";
defparam \E_ctrl_invalidate_i~0 .lut_mask = 64'h9669699696696996;
defparam \E_ctrl_invalidate_i~0 .shared_arith = "off";

cyclonev_lcell_comb \E_ctrl_invalidate_i~1 (
	.dataa(!\E_iw[14]~q ),
	.datab(!\Equal239~0_combout ),
	.datac(!\E_ctrl_invalidate_i~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_ctrl_invalidate_i~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_ctrl_invalidate_i~1 .extended_lut = "off";
defparam \E_ctrl_invalidate_i~1 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \E_ctrl_invalidate_i~1 .shared_arith = "off";

dffeas M_ctrl_invalidate_i(
	.clk(clk_clk),
	.d(\E_ctrl_invalidate_i~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_ctrl_invalidate_i~q ),
	.prn(vcc));
defparam M_ctrl_invalidate_i.is_wysiwyg = "true";
defparam M_ctrl_invalidate_i.power_up = "low";

dffeas A_ctrl_invalidate_i(
	.clk(clk_clk),
	.d(\M_ctrl_invalidate_i~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\A_ctrl_invalidate_i~q ),
	.prn(vcc));
defparam A_ctrl_invalidate_i.is_wysiwyg = "true";
defparam A_ctrl_invalidate_i.power_up = "low";

cyclonev_lcell_comb ic_fill_prevent_refill_nxt(
	.dataa(!\A_valid_from_M~q ),
	.datab(!\ic_fill_prevent_refill~q ),
	.datac(!\D_ic_fill_starting~combout ),
	.datad(!\A_ctrl_invalidate_i~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_prevent_refill_nxt~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam ic_fill_prevent_refill_nxt.extended_lut = "off";
defparam ic_fill_prevent_refill_nxt.lut_mask = 64'hFFBFFFBFFFBFFFBF;
defparam ic_fill_prevent_refill_nxt.shared_arith = "off";

dffeas ic_fill_prevent_refill(
	.clk(clk_clk),
	.d(\ic_fill_prevent_refill_nxt~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ic_fill_prevent_refill~q ),
	.prn(vcc));
defparam ic_fill_prevent_refill.is_wysiwyg = "true";
defparam ic_fill_prevent_refill.power_up = "low";

cyclonev_lcell_comb \D_ic_fill_starting~0 (
	.dataa(!\D_ic_fill_same_tag_line~q ),
	.datab(!\ic_fill_prevent_refill~q ),
	.datac(!\ic_fill_active~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ic_fill_starting~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ic_fill_starting~0 .extended_lut = "off";
defparam \D_ic_fill_starting~0 .lut_mask = 64'hFEFEFEFEFEFEFEFE;
defparam \D_ic_fill_starting~0 .shared_arith = "off";

cyclonev_lcell_comb D_ic_fill_starting(
	.dataa(!\M_pipe_flush~q ),
	.datab(!\E_valid_jmp_indirect~q ),
	.datac(!\D_iw_valid~q ),
	.datad(!\D_kill~q ),
	.datae(!\D_ic_fill_starting~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ic_fill_starting~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam D_ic_fill_starting.extended_lut = "off";
defparam D_ic_fill_starting.lut_mask = 64'hFFFDFFFFFFFDFFFF;
defparam D_ic_fill_starting.shared_arith = "off";

dffeas \ic_fill_initial_offset[2] (
	.clk(clk_clk),
	.d(\D_pc[2]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\D_ic_fill_starting~combout ),
	.q(\ic_fill_initial_offset[2]~q ),
	.prn(vcc));
defparam \ic_fill_initial_offset[2] .is_wysiwyg = "true";
defparam \ic_fill_initial_offset[2] .power_up = "low";

dffeas D_ic_fill_starting_d1(
	.clk(clk_clk),
	.d(\D_ic_fill_starting~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\D_ic_fill_starting_d1~q ),
	.prn(vcc));
defparam D_ic_fill_starting_d1.is_wysiwyg = "true";
defparam D_ic_fill_starting_d1.power_up = "low";

dffeas \ic_fill_initial_offset[0] (
	.clk(clk_clk),
	.d(\D_pc[0]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\D_ic_fill_starting~combout ),
	.q(\ic_fill_initial_offset[0]~q ),
	.prn(vcc));
defparam \ic_fill_initial_offset[0] .is_wysiwyg = "true";
defparam \ic_fill_initial_offset[0] .power_up = "low";

cyclonev_lcell_comb \ic_fill_dp_offset_nxt[0]~1 (
	.dataa(!\ic_fill_initial_offset[0]~q ),
	.datab(!\D_ic_fill_starting_d1~q ),
	.datac(!\ic_fill_dp_offset[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_dp_offset_nxt[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_dp_offset_nxt[0]~1 .extended_lut = "off";
defparam \ic_fill_dp_offset_nxt[0]~1 .lut_mask = 64'hD1D1D1D1D1D1D1D1;
defparam \ic_fill_dp_offset_nxt[0]~1 .shared_arith = "off";

dffeas i_readdatavalid_d1(
	.clk(clk_clk),
	.d(WideOr15),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdatavalid_d1~q ),
	.prn(vcc));
defparam i_readdatavalid_d1.is_wysiwyg = "true";
defparam i_readdatavalid_d1.power_up = "low";

cyclonev_lcell_comb \ic_fill_dp_offset_en~0 (
	.dataa(!\i_readdatavalid_d1~q ),
	.datab(!\D_ic_fill_starting_d1~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_dp_offset_en~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_dp_offset_en~0 .extended_lut = "off";
defparam \ic_fill_dp_offset_en~0 .lut_mask = 64'h7777777777777777;
defparam \ic_fill_dp_offset_en~0 .shared_arith = "off";

dffeas \ic_fill_dp_offset[0] (
	.clk(clk_clk),
	.d(\ic_fill_dp_offset_nxt[0]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ic_fill_dp_offset_en~0_combout ),
	.q(\ic_fill_dp_offset[0]~q ),
	.prn(vcc));
defparam \ic_fill_dp_offset[0] .is_wysiwyg = "true";
defparam \ic_fill_dp_offset[0] .power_up = "low";

dffeas \ic_fill_initial_offset[1] (
	.clk(clk_clk),
	.d(\D_pc[1]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\D_ic_fill_starting~combout ),
	.q(\ic_fill_initial_offset[1]~q ),
	.prn(vcc));
defparam \ic_fill_initial_offset[1] .is_wysiwyg = "true";
defparam \ic_fill_initial_offset[1] .power_up = "low";

cyclonev_lcell_comb \ic_fill_dp_offset_nxt[1]~2 (
	.dataa(!\D_ic_fill_starting_d1~q ),
	.datab(!\ic_fill_dp_offset[0]~q ),
	.datac(!\ic_fill_initial_offset[1]~q ),
	.datad(!\ic_fill_dp_offset[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_dp_offset_nxt[1]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_dp_offset_nxt[1]~2 .extended_lut = "off";
defparam \ic_fill_dp_offset_nxt[1]~2 .lut_mask = 64'h9F6F9F6F9F6F9F6F;
defparam \ic_fill_dp_offset_nxt[1]~2 .shared_arith = "off";

dffeas \ic_fill_dp_offset[1] (
	.clk(clk_clk),
	.d(\ic_fill_dp_offset_nxt[1]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ic_fill_dp_offset_en~0_combout ),
	.q(\ic_fill_dp_offset[1]~q ),
	.prn(vcc));
defparam \ic_fill_dp_offset[1] .is_wysiwyg = "true";
defparam \ic_fill_dp_offset[1] .power_up = "low";

dffeas \ic_fill_dp_offset[2] (
	.clk(clk_clk),
	.d(\ic_fill_dp_offset_nxt[2]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ic_fill_dp_offset_en~0_combout ),
	.q(\ic_fill_dp_offset[2]~q ),
	.prn(vcc));
defparam \ic_fill_dp_offset[2] .is_wysiwyg = "true";
defparam \ic_fill_dp_offset[2] .power_up = "low";

cyclonev_lcell_comb \ic_fill_dp_offset_nxt[2]~0 (
	.dataa(!\D_ic_fill_starting_d1~q ),
	.datab(!\ic_fill_dp_offset[0]~q ),
	.datac(!\ic_fill_dp_offset[1]~q ),
	.datad(!\ic_fill_initial_offset[2]~q ),
	.datae(!\ic_fill_dp_offset[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_dp_offset_nxt[2]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_dp_offset_nxt[2]~0 .extended_lut = "off";
defparam \ic_fill_dp_offset_nxt[2]~0 .lut_mask = 64'h69FF96FF69FF96FF;
defparam \ic_fill_dp_offset_nxt[2]~0 .shared_arith = "off";

cyclonev_lcell_comb \ic_fill_active_nxt~0 (
	.dataa(!\i_readdatavalid_d1~q ),
	.datab(!\ic_fill_initial_offset[0]~q ),
	.datac(!\ic_fill_dp_offset_nxt[0]~1_combout ),
	.datad(!\ic_fill_initial_offset[1]~q ),
	.datae(!\ic_fill_dp_offset_nxt[1]~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_active_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_active_nxt~0 .extended_lut = "off";
defparam \ic_fill_active_nxt~0 .lut_mask = 64'h7DD7D77D7DD7D77D;
defparam \ic_fill_active_nxt~0 .shared_arith = "off";

cyclonev_lcell_comb \ic_fill_active_nxt~1 (
	.dataa(!\ic_fill_active~q ),
	.datab(!\D_ic_fill_starting~combout ),
	.datac(!\ic_fill_initial_offset[2]~q ),
	.datad(!\ic_fill_dp_offset_nxt[2]~0_combout ),
	.datae(!\ic_fill_active_nxt~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_active_nxt~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_active_nxt~1 .extended_lut = "off";
defparam \ic_fill_active_nxt~1 .lut_mask = 64'hFFFF7FF7FFFF7FF7;
defparam \ic_fill_active_nxt~1 .shared_arith = "off";

dffeas ic_fill_active(
	.clk(clk_clk),
	.d(\ic_fill_active_nxt~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ic_fill_active~q ),
	.prn(vcc));
defparam ic_fill_active.is_wysiwyg = "true";
defparam ic_fill_active.power_up = "low";

cyclonev_lcell_comb \ic_fill_ap_cnt_nxt[0]~3 (
	.dataa(!nonposted_cmd_accepted),
	.datab(!\ic_fill_ap_cnt[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_ap_cnt_nxt[0]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_ap_cnt_nxt[0]~3 .extended_lut = "off";
defparam \ic_fill_ap_cnt_nxt[0]~3 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \ic_fill_ap_cnt_nxt[0]~3 .shared_arith = "off";

cyclonev_lcell_comb \ic_fill_ap_offset[2]~0 (
	.dataa(!save_dest_id),
	.datab(!WideOr0),
	.datac(!\D_ic_fill_starting~combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_ap_offset[2]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_ap_offset[2]~0 .extended_lut = "off";
defparam \ic_fill_ap_offset[2]~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \ic_fill_ap_offset[2]~0 .shared_arith = "off";

dffeas \ic_fill_ap_cnt[0] (
	.clk(clk_clk),
	.d(\ic_fill_ap_cnt_nxt[0]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ic_fill_ap_offset[2]~0_combout ),
	.q(\ic_fill_ap_cnt[0]~q ),
	.prn(vcc));
defparam \ic_fill_ap_cnt[0] .is_wysiwyg = "true";
defparam \ic_fill_ap_cnt[0] .power_up = "low";

cyclonev_lcell_comb \ic_fill_ap_cnt_nxt[1]~2 (
	.dataa(!nonposted_cmd_accepted),
	.datab(!\ic_fill_ap_cnt[1]~q ),
	.datac(!\ic_fill_ap_cnt[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_ap_cnt_nxt[1]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_ap_cnt_nxt[1]~2 .extended_lut = "off";
defparam \ic_fill_ap_cnt_nxt[1]~2 .lut_mask = 64'h7D7D7D7D7D7D7D7D;
defparam \ic_fill_ap_cnt_nxt[1]~2 .shared_arith = "off";

dffeas \ic_fill_ap_cnt[1] (
	.clk(clk_clk),
	.d(\ic_fill_ap_cnt_nxt[1]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ic_fill_ap_offset[2]~0_combout ),
	.q(\ic_fill_ap_cnt[1]~q ),
	.prn(vcc));
defparam \ic_fill_ap_cnt[1] .is_wysiwyg = "true";
defparam \ic_fill_ap_cnt[1] .power_up = "low";

cyclonev_lcell_comb \ic_fill_ap_cnt_nxt[2]~1 (
	.dataa(!nonposted_cmd_accepted),
	.datab(!\ic_fill_ap_cnt[2]~q ),
	.datac(!\ic_fill_ap_cnt[1]~q ),
	.datad(!\ic_fill_ap_cnt[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_ap_cnt_nxt[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_ap_cnt_nxt[2]~1 .extended_lut = "off";
defparam \ic_fill_ap_cnt_nxt[2]~1 .lut_mask = 64'hD77DD77DD77DD77D;
defparam \ic_fill_ap_cnt_nxt[2]~1 .shared_arith = "off";

dffeas \ic_fill_ap_cnt[2] (
	.clk(clk_clk),
	.d(\ic_fill_ap_cnt_nxt[2]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ic_fill_ap_offset[2]~0_combout ),
	.q(\ic_fill_ap_cnt[2]~q ),
	.prn(vcc));
defparam \ic_fill_ap_cnt[2] .is_wysiwyg = "true";
defparam \ic_fill_ap_cnt[2] .power_up = "low";

cyclonev_lcell_comb \ic_fill_ap_cnt_nxt[3]~0 (
	.dataa(!nonposted_cmd_accepted),
	.datab(!\ic_fill_ap_cnt[3]~q ),
	.datac(!\ic_fill_ap_cnt[2]~q ),
	.datad(!\ic_fill_ap_cnt[1]~q ),
	.datae(!\ic_fill_ap_cnt[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_ap_cnt_nxt[3]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_ap_cnt_nxt[3]~0 .extended_lut = "off";
defparam \ic_fill_ap_cnt_nxt[3]~0 .lut_mask = 64'h7DD7D77D7DD7D77D;
defparam \ic_fill_ap_cnt_nxt[3]~0 .shared_arith = "off";

dffeas \ic_fill_ap_cnt[3] (
	.clk(clk_clk),
	.d(\ic_fill_ap_cnt_nxt[3]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ic_fill_ap_offset[2]~0_combout ),
	.q(\ic_fill_ap_cnt[3]~q ),
	.prn(vcc));
defparam \ic_fill_ap_cnt[3] .is_wysiwyg = "true";
defparam \ic_fill_ap_cnt[3] .power_up = "low";

cyclonev_lcell_comb \i_read_nxt~0 (
	.dataa(!clr_break_line1),
	.datab(!\ic_fill_active~q ),
	.datac(!\ic_fill_ap_cnt[3]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\i_read_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \i_read_nxt~0 .extended_lut = "off";
defparam \i_read_nxt~0 .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \i_read_nxt~0 .shared_arith = "off";

cyclonev_lcell_comb \i_read_nxt~1 (
	.dataa(!i_read1),
	.datab(!suppress_change_dest_id),
	.datac(!WideOr0),
	.datad(!\i_read_nxt~0_combout ),
	.datae(!\D_ic_fill_starting~combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\i_read_nxt~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \i_read_nxt~1 .extended_lut = "off";
defparam \i_read_nxt~1 .lut_mask = 64'hFFF7FFFFFFF7FFFF;
defparam \i_read_nxt~1 .shared_arith = "off";

cyclonev_lcell_comb \ic_fill_ap_offset_nxt[0]~0 (
	.dataa(!ic_fill_ap_offset_0),
	.datab(!nonposted_cmd_accepted),
	.datac(!\D_pc[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_ap_offset_nxt[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_ap_offset_nxt[0]~0 .extended_lut = "off";
defparam \ic_fill_ap_offset_nxt[0]~0 .lut_mask = 64'h8B8B8B8B8B8B8B8B;
defparam \ic_fill_ap_offset_nxt[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \ic_tag_wraddress_nxt~0 (
	.dataa(!ic_fill_line_0),
	.datab(!\D_ic_fill_starting~combout ),
	.datac(!\D_pc[3]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_tag_wraddress_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_tag_wraddress_nxt~0 .extended_lut = "off";
defparam \ic_tag_wraddress_nxt~0 .lut_mask = 64'h4747474747474747;
defparam \ic_tag_wraddress_nxt~0 .shared_arith = "off";

cyclonev_lcell_comb \ic_fill_ap_offset_nxt[2]~1 (
	.dataa(!ic_fill_ap_offset_0),
	.datab(!ic_fill_ap_offset_2),
	.datac(!ic_fill_ap_offset_1),
	.datad(!nonposted_cmd_accepted),
	.datae(!\D_pc[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_ap_offset_nxt[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_ap_offset_nxt[2]~1 .extended_lut = "off";
defparam \ic_fill_ap_offset_nxt[2]~1 .lut_mask = 64'h6996FFFF6996FFFF;
defparam \ic_fill_ap_offset_nxt[2]~1 .shared_arith = "off";

cyclonev_lcell_comb \ic_fill_ap_offset_nxt[1]~2 (
	.dataa(!ic_fill_ap_offset_0),
	.datab(!ic_fill_ap_offset_1),
	.datac(!nonposted_cmd_accepted),
	.datad(!\D_pc[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_ap_offset_nxt[1]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_ap_offset_nxt[1]~2 .extended_lut = "off";
defparam \ic_fill_ap_offset_nxt[1]~2 .lut_mask = 64'h96FF96FF96FF96FF;
defparam \ic_fill_ap_offset_nxt[1]~2 .shared_arith = "off";

cyclonev_lcell_comb \ic_tag_wraddress_nxt~1 (
	.dataa(!ic_fill_line_5),
	.datab(!\D_ic_fill_starting~combout ),
	.datac(!\D_pc[8]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_tag_wraddress_nxt~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_tag_wraddress_nxt~1 .extended_lut = "off";
defparam \ic_tag_wraddress_nxt~1 .lut_mask = 64'h4747474747474747;
defparam \ic_tag_wraddress_nxt~1 .shared_arith = "off";

cyclonev_lcell_comb \ic_tag_wraddress_nxt~2 (
	.dataa(!ic_fill_line_4),
	.datab(!\D_ic_fill_starting~combout ),
	.datac(!\D_pc[7]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_tag_wraddress_nxt~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_tag_wraddress_nxt~2 .extended_lut = "off";
defparam \ic_tag_wraddress_nxt~2 .lut_mask = 64'h4747474747474747;
defparam \ic_tag_wraddress_nxt~2 .shared_arith = "off";

cyclonev_lcell_comb \ic_tag_wraddress_nxt~3 (
	.dataa(!ic_fill_line_3),
	.datab(!\D_ic_fill_starting~combout ),
	.datac(!\D_pc[6]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_tag_wraddress_nxt~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_tag_wraddress_nxt~3 .extended_lut = "off";
defparam \ic_tag_wraddress_nxt~3 .lut_mask = 64'h4747474747474747;
defparam \ic_tag_wraddress_nxt~3 .shared_arith = "off";

cyclonev_lcell_comb \ic_tag_wraddress_nxt~4 (
	.dataa(!ic_fill_line_2),
	.datab(!\D_ic_fill_starting~combout ),
	.datac(!\D_pc[5]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_tag_wraddress_nxt~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_tag_wraddress_nxt~4 .extended_lut = "off";
defparam \ic_tag_wraddress_nxt~4 .lut_mask = 64'h4747474747474747;
defparam \ic_tag_wraddress_nxt~4 .shared_arith = "off";

cyclonev_lcell_comb \ic_tag_wraddress_nxt~5 (
	.dataa(!ic_fill_line_1),
	.datab(!\D_ic_fill_starting~combout ),
	.datac(!\D_pc[4]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_tag_wraddress_nxt~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_tag_wraddress_nxt~5 .extended_lut = "off";
defparam \ic_tag_wraddress_nxt~5 .lut_mask = 64'h4747474747474747;
defparam \ic_tag_wraddress_nxt~5 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_mem16~0 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[3]~q ),
	.datac(!\D_iw[4]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_mem16~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_mem16~0 .extended_lut = "off";
defparam \D_ctrl_mem16~0 .lut_mask = 64'hF7F7F7F7F7F7F7F7;
defparam \D_ctrl_mem16~0 .shared_arith = "off";

dffeas E_ctrl_mem16(
	.clk(clk_clk),
	.d(\D_ctrl_mem16~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_ctrl_mem16~q ),
	.prn(vcc));
defparam E_ctrl_mem16.is_wysiwyg = "true";
defparam E_ctrl_mem16.power_up = "low";

cyclonev_lcell_comb \D_ctrl_mem8~0 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[1]~q ),
	.datac(!\D_iw[2]~q ),
	.datad(!\D_iw[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_mem8~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_mem8~0 .extended_lut = "off";
defparam \D_ctrl_mem8~0 .lut_mask = 64'hFF7FFF7FFF7FFF7F;
defparam \D_ctrl_mem8~0 .shared_arith = "off";

dffeas E_ctrl_mem8(
	.clk(clk_clk),
	.d(\D_ctrl_mem8~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\D_iw[4]~q ),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_ctrl_mem8~q ),
	.prn(vcc));
defparam E_ctrl_mem8.is_wysiwyg = "true";
defparam E_ctrl_mem8.power_up = "low";

cyclonev_lcell_comb \E_mem_byte_en~0 (
	.dataa(!\Add9~65_sumout ),
	.datab(!\Add9~69_sumout ),
	.datac(!\E_ctrl_mem16~q ),
	.datad(!\E_ctrl_mem8~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_mem_byte_en~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_mem_byte_en~0 .extended_lut = "off";
defparam \E_mem_byte_en~0 .lut_mask = 64'hEFFEEFFEEFFEEFFE;
defparam \E_mem_byte_en~0 .shared_arith = "off";

dffeas \M_mem_byte_en[0] (
	.clk(clk_clk),
	.d(\E_mem_byte_en~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_mem_byte_en[0]~q ),
	.prn(vcc));
defparam \M_mem_byte_en[0] .is_wysiwyg = "true";
defparam \M_mem_byte_en[0] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[16]~73 (
	.dataa(!\D_src2_reg[0]~4_combout ),
	.datab(!\D_src2_reg[0]~5_combout ),
	.datac(!\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[16] ),
	.datad(!\E_alu_result[16]~combout ),
	.datae(!\D_src2_reg[16]~61_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[16]~73_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[16]~73 .extended_lut = "off";
defparam \D_src2_reg[16]~73 .lut_mask = 64'h47FFFFFF47FFFFFF;
defparam \D_src2_reg[16]~73 .shared_arith = "off";

dffeas \E_src2_reg[16] (
	.clk(clk_clk),
	.d(\D_src2_reg[16]~73_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_src2_reg[16]~q ),
	.prn(vcc));
defparam \E_src2_reg[16] .is_wysiwyg = "true";
defparam \E_src2_reg[16] .power_up = "low";

cyclonev_lcell_comb \E_st_data[23]~0 (
	.dataa(!\E_ctrl_mem16~q ),
	.datab(!\E_ctrl_mem8~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_st_data[23]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_st_data[23]~0 .extended_lut = "off";
defparam \E_st_data[23]~0 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \E_st_data[23]~0 .shared_arith = "off";

dffeas \M_st_data[16] (
	.clk(clk_clk),
	.d(\E_src2_reg[0]~q ),
	.asdata(\E_src2_reg[16]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_st_data[23]~0_combout ),
	.ena(!\A_mem_stall~q ),
	.q(\M_st_data[16]~q ),
	.prn(vcc));
defparam \M_st_data[16] .is_wysiwyg = "true";
defparam \M_st_data[16] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[22]~74 (
	.dataa(!\D_src2_reg[0]~4_combout ),
	.datab(!\D_src2_reg[0]~5_combout ),
	.datac(!\E_alu_result[22]~combout ),
	.datad(!\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[22] ),
	.datae(!\D_src2_reg[22]~26_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[22]~74_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[22]~74 .extended_lut = "off";
defparam \D_src2_reg[22]~74 .lut_mask = 64'h47FFFFFF47FFFFFF;
defparam \D_src2_reg[22]~74 .shared_arith = "off";

dffeas \E_src2_reg[22] (
	.clk(clk_clk),
	.d(\D_src2_reg[22]~74_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_src2_reg[22]~q ),
	.prn(vcc));
defparam \E_src2_reg[22] .is_wysiwyg = "true";
defparam \E_src2_reg[22] .power_up = "low";

dffeas \M_st_data[22] (
	.clk(clk_clk),
	.d(\E_src2_reg[6]~q ),
	.asdata(\E_src2_reg[22]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_st_data[23]~0_combout ),
	.ena(!\A_mem_stall~q ),
	.q(\M_st_data[22]~q ),
	.prn(vcc));
defparam \M_st_data[22] .is_wysiwyg = "true";
defparam \M_st_data[22] .power_up = "low";

cyclonev_lcell_comb \E_mem_byte_en[2]~1 (
	.dataa(!\Add9~65_sumout ),
	.datab(!\Add9~69_sumout ),
	.datac(!\E_ctrl_mem16~q ),
	.datad(!\E_ctrl_mem8~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_mem_byte_en[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_mem_byte_en[2]~1 .extended_lut = "off";
defparam \E_mem_byte_en[2]~1 .lut_mask = 64'hBFFBBFFBBFFBBFFB;
defparam \E_mem_byte_en[2]~1 .shared_arith = "off";

dffeas \M_mem_byte_en[2] (
	.clk(clk_clk),
	.d(\E_mem_byte_en[2]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_mem_byte_en[2]~q ),
	.prn(vcc));
defparam \M_mem_byte_en[2] .is_wysiwyg = "true";
defparam \M_mem_byte_en[2] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[23]~75 (
	.dataa(!\D_src2_reg[23]~28_combout ),
	.datab(!\Equal304~0_combout ),
	.datac(!\D_src2_reg[0]~0_combout ),
	.datad(!\D_src2_reg[0]~1_combout ),
	.datae(!\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[23] ),
	.dataf(!\D_src2_reg[23]~27_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[23]~75_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[23]~75 .extended_lut = "off";
defparam \D_src2_reg[23]~75 .lut_mask = 64'hFFFDFFFFFFFFFFFF;
defparam \D_src2_reg[23]~75 .shared_arith = "off";

dffeas \E_src2_reg[23] (
	.clk(clk_clk),
	.d(\D_src2_reg[23]~75_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_src2_reg[23]~q ),
	.prn(vcc));
defparam \E_src2_reg[23] .is_wysiwyg = "true";
defparam \E_src2_reg[23] .power_up = "low";

dffeas \M_st_data[23] (
	.clk(clk_clk),
	.d(\E_src2_reg[7]~q ),
	.asdata(\E_src2_reg[23]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_st_data[23]~0_combout ),
	.ena(!\A_mem_stall~q ),
	.q(\M_st_data[23]~q ),
	.prn(vcc));
defparam \M_st_data[23] .is_wysiwyg = "true";
defparam \M_st_data[23] .power_up = "low";

dffeas \E_src2_reg[8] (
	.clk(clk_clk),
	.d(\D_src2_reg[8]~49_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_src2_reg[8]~q ),
	.prn(vcc));
defparam \E_src2_reg[8] .is_wysiwyg = "true";
defparam \E_src2_reg[8] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[24]~76 (
	.dataa(!\D_src2_reg[24]~30_combout ),
	.datab(!\Equal304~0_combout ),
	.datac(!\D_src2_reg[0]~0_combout ),
	.datad(!\D_src2_reg[0]~1_combout ),
	.datae(!\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[24] ),
	.dataf(!\D_src2_reg[24]~29_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[24]~76_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[24]~76 .extended_lut = "off";
defparam \D_src2_reg[24]~76 .lut_mask = 64'hFFFDFFFFFFFFFFFF;
defparam \D_src2_reg[24]~76 .shared_arith = "off";

dffeas \E_src2_reg[24] (
	.clk(clk_clk),
	.d(\D_src2_reg[24]~76_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_src2_reg[24]~q ),
	.prn(vcc));
defparam \E_src2_reg[24] .is_wysiwyg = "true";
defparam \E_src2_reg[24] .power_up = "low";

cyclonev_lcell_comb \E_st_data[24]~1 (
	.dataa(!\E_ctrl_mem16~q ),
	.datab(!\E_src2_reg[8]~q ),
	.datac(!\E_src2_reg[24]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_st_data[24]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_st_data[24]~1 .extended_lut = "off";
defparam \E_st_data[24]~1 .lut_mask = 64'h2727272727272727;
defparam \E_st_data[24]~1 .shared_arith = "off";

dffeas \M_st_data[24] (
	.clk(clk_clk),
	.d(\E_st_data[24]~1_combout ),
	.asdata(\E_src2_reg[0]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_ctrl_mem8~q ),
	.ena(!\A_mem_stall~q ),
	.q(\M_st_data[24]~q ),
	.prn(vcc));
defparam \M_st_data[24] .is_wysiwyg = "true";
defparam \M_st_data[24] .power_up = "low";

cyclonev_lcell_comb \E_mem_byte_en[3]~2 (
	.dataa(!\Add9~65_sumout ),
	.datab(!\Add9~69_sumout ),
	.datac(!\E_ctrl_mem16~q ),
	.datad(!\E_ctrl_mem8~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_mem_byte_en[3]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_mem_byte_en[3]~2 .extended_lut = "off";
defparam \E_mem_byte_en[3]~2 .lut_mask = 64'h7FF77FF77FF77FF7;
defparam \E_mem_byte_en[3]~2 .shared_arith = "off";

dffeas \M_mem_byte_en[3] (
	.clk(clk_clk),
	.d(\E_mem_byte_en[3]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_mem_byte_en[3]~q ),
	.prn(vcc));
defparam \M_mem_byte_en[3] .is_wysiwyg = "true";
defparam \M_mem_byte_en[3] .power_up = "low";

dffeas \E_src2_reg[9] (
	.clk(clk_clk),
	.d(\D_src2_reg[9]~51_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_src2_reg[9]~q ),
	.prn(vcc));
defparam \E_src2_reg[9] .is_wysiwyg = "true";
defparam \E_src2_reg[9] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[25]~77 (
	.dataa(!\D_src2_reg[25]~32_combout ),
	.datab(!\Equal304~0_combout ),
	.datac(!\D_src2_reg[0]~0_combout ),
	.datad(!\D_src2_reg[0]~1_combout ),
	.datae(!\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[25] ),
	.dataf(!\D_src2_reg[25]~31_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[25]~77_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[25]~77 .extended_lut = "off";
defparam \D_src2_reg[25]~77 .lut_mask = 64'hFFFDFFFFFFFFFFFF;
defparam \D_src2_reg[25]~77 .shared_arith = "off";

dffeas \E_src2_reg[25] (
	.clk(clk_clk),
	.d(\D_src2_reg[25]~77_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_src2_reg[25]~q ),
	.prn(vcc));
defparam \E_src2_reg[25] .is_wysiwyg = "true";
defparam \E_src2_reg[25] .power_up = "low";

cyclonev_lcell_comb \E_st_data[25]~2 (
	.dataa(!\E_ctrl_mem16~q ),
	.datab(!\E_src2_reg[9]~q ),
	.datac(!\E_src2_reg[25]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_st_data[25]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_st_data[25]~2 .extended_lut = "off";
defparam \E_st_data[25]~2 .lut_mask = 64'h2727272727272727;
defparam \E_st_data[25]~2 .shared_arith = "off";

dffeas \M_st_data[25] (
	.clk(clk_clk),
	.d(\E_st_data[25]~2_combout ),
	.asdata(\E_src2_reg[1]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_ctrl_mem8~q ),
	.ena(!\A_mem_stall~q ),
	.q(\M_st_data[25]~q ),
	.prn(vcc));
defparam \M_st_data[25] .is_wysiwyg = "true";
defparam \M_st_data[25] .power_up = "low";

dffeas \E_src2_reg[15] (
	.clk(clk_clk),
	.d(\D_src2_reg[15]~63_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_src2_reg[15]~q ),
	.prn(vcc));
defparam \E_src2_reg[15] .is_wysiwyg = "true";
defparam \E_src2_reg[15] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[31]~89 (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\Add9~73_sumout ),
	.datac(!\E_alu_result~10_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[31]~89_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[31]~89 .extended_lut = "off";
defparam \D_src2_reg[31]~89 .lut_mask = 64'hFEFEFEFEFEFEFEFE;
defparam \D_src2_reg[31]~89 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[31]~78 (
	.dataa(!\D_src2_reg[0]~2_combout ),
	.datab(!\D_src2_reg[31]~36_combout ),
	.datac(!\D_src2_reg[0]~4_combout ),
	.datad(!\D_src2_reg[0]~5_combout ),
	.datae(!\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[31] ),
	.dataf(!\D_src2_reg[31]~89_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[31]~78_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[31]~78 .extended_lut = "off";
defparam \D_src2_reg[31]~78 .lut_mask = 64'hFFFFFFFFFF7FFFFF;
defparam \D_src2_reg[31]~78 .shared_arith = "off";

dffeas \E_src2_reg[31] (
	.clk(clk_clk),
	.d(\D_src2_reg[31]~78_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_src2_reg[31]~q ),
	.prn(vcc));
defparam \E_src2_reg[31] .is_wysiwyg = "true";
defparam \E_src2_reg[31] .power_up = "low";

cyclonev_lcell_comb \E_st_data[31]~3 (
	.dataa(!\E_ctrl_mem16~q ),
	.datab(!\E_src2_reg[15]~q ),
	.datac(!\E_src2_reg[31]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_st_data[31]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_st_data[31]~3 .extended_lut = "off";
defparam \E_st_data[31]~3 .lut_mask = 64'h2727272727272727;
defparam \E_st_data[31]~3 .shared_arith = "off";

dffeas \M_st_data[31] (
	.clk(clk_clk),
	.d(\E_st_data[31]~3_combout ),
	.asdata(\E_src2_reg[7]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_ctrl_mem8~q ),
	.ena(!\A_mem_stall~q ),
	.q(\M_st_data[31]~q ),
	.prn(vcc));
defparam \M_st_data[31] .is_wysiwyg = "true";
defparam \M_st_data[31] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[21]~79 (
	.dataa(!\D_src2_reg[0]~4_combout ),
	.datab(!\D_src2_reg[0]~5_combout ),
	.datac(!\E_alu_result[21]~combout ),
	.datad(!\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[21] ),
	.datae(!\D_src2_reg[21]~37_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[21]~79_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[21]~79 .extended_lut = "off";
defparam \D_src2_reg[21]~79 .lut_mask = 64'h47FFFFFF47FFFFFF;
defparam \D_src2_reg[21]~79 .shared_arith = "off";

dffeas \E_src2_reg[21] (
	.clk(clk_clk),
	.d(\D_src2_reg[21]~79_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_src2_reg[21]~q ),
	.prn(vcc));
defparam \E_src2_reg[21] .is_wysiwyg = "true";
defparam \E_src2_reg[21] .power_up = "low";

dffeas \M_st_data[21] (
	.clk(clk_clk),
	.d(\E_src2_reg[5]~q ),
	.asdata(\E_src2_reg[21]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_st_data[23]~0_combout ),
	.ena(!\A_mem_stall~q ),
	.q(\M_st_data[21]~q ),
	.prn(vcc));
defparam \M_st_data[21] .is_wysiwyg = "true";
defparam \M_st_data[21] .power_up = "low";

dffeas \E_src2_reg[11] (
	.clk(clk_clk),
	.d(\D_src2_reg[11]~39_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_src2_reg[11]~q ),
	.prn(vcc));
defparam \E_src2_reg[11] .is_wysiwyg = "true";
defparam \E_src2_reg[11] .power_up = "low";

dffeas \M_st_data[11] (
	.clk(clk_clk),
	.d(\E_src2_reg[3]~q ),
	.asdata(\E_src2_reg[11]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\E_ctrl_mem8~q ),
	.ena(!\A_mem_stall~q ),
	.q(\M_st_data[11]~q ),
	.prn(vcc));
defparam \M_st_data[11] .is_wysiwyg = "true";
defparam \M_st_data[11] .power_up = "low";

cyclonev_lcell_comb \E_mem_byte_en[1]~3 (
	.dataa(!\Add9~65_sumout ),
	.datab(!\Add9~69_sumout ),
	.datac(!\E_ctrl_mem16~q ),
	.datad(!\E_ctrl_mem8~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_mem_byte_en[1]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_mem_byte_en[1]~3 .extended_lut = "off";
defparam \E_mem_byte_en[1]~3 .lut_mask = 64'hDFFDDFFDDFFDDFFD;
defparam \E_mem_byte_en[1]~3 .shared_arith = "off";

dffeas \M_mem_byte_en[1] (
	.clk(clk_clk),
	.d(\E_mem_byte_en[1]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\M_mem_byte_en[1]~q ),
	.prn(vcc));
defparam \M_mem_byte_en[1] .is_wysiwyg = "true";
defparam \M_mem_byte_en[1] .power_up = "low";

dffeas \E_src2_reg[12] (
	.clk(clk_clk),
	.d(\D_src2_reg[12]~65_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_src2_reg[12]~q ),
	.prn(vcc));
defparam \E_src2_reg[12] .is_wysiwyg = "true";
defparam \E_src2_reg[12] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[28]~80 (
	.dataa(!\D_src2_reg[28]~42_combout ),
	.datab(!\Equal304~0_combout ),
	.datac(!\D_src2_reg[0]~0_combout ),
	.datad(!\D_src2_reg[0]~1_combout ),
	.datae(!\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[28] ),
	.dataf(!\D_src2_reg[28]~40_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[28]~80_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[28]~80 .extended_lut = "off";
defparam \D_src2_reg[28]~80 .lut_mask = 64'hFFFDFFFFFFFFFFFF;
defparam \D_src2_reg[28]~80 .shared_arith = "off";

dffeas \E_src2_reg[28] (
	.clk(clk_clk),
	.d(\D_src2_reg[28]~80_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_src2_reg[28]~q ),
	.prn(vcc));
defparam \E_src2_reg[28] .is_wysiwyg = "true";
defparam \E_src2_reg[28] .power_up = "low";

cyclonev_lcell_comb \E_st_data[28]~4 (
	.dataa(!\E_ctrl_mem16~q ),
	.datab(!\E_src2_reg[12]~q ),
	.datac(!\E_src2_reg[28]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_st_data[28]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_st_data[28]~4 .extended_lut = "off";
defparam \E_st_data[28]~4 .lut_mask = 64'h2727272727272727;
defparam \E_st_data[28]~4 .shared_arith = "off";

dffeas \M_st_data[28] (
	.clk(clk_clk),
	.d(\E_st_data[28]~4_combout ),
	.asdata(\E_src2_reg[4]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_ctrl_mem8~q ),
	.ena(!\A_mem_stall~q ),
	.q(\M_st_data[28]~q ),
	.prn(vcc));
defparam \M_st_data[28] .is_wysiwyg = "true";
defparam \M_st_data[28] .power_up = "low";

dffeas \E_src2_reg[10] (
	.clk(clk_clk),
	.d(\D_src2_reg[10]~44_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_src2_reg[10]~q ),
	.prn(vcc));
defparam \E_src2_reg[10] .is_wysiwyg = "true";
defparam \E_src2_reg[10] .power_up = "low";

dffeas \M_st_data[10] (
	.clk(clk_clk),
	.d(\E_src2_reg[2]~q ),
	.asdata(\E_src2_reg[10]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\E_ctrl_mem8~q ),
	.ena(!\A_mem_stall~q ),
	.q(\M_st_data[10]~q ),
	.prn(vcc));
defparam \M_st_data[10] .is_wysiwyg = "true";
defparam \M_st_data[10] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[27]~81 (
	.dataa(!\D_src2_reg[27]~47_combout ),
	.datab(!\Equal304~0_combout ),
	.datac(!\D_src2_reg[0]~0_combout ),
	.datad(!\D_src2_reg[0]~1_combout ),
	.datae(!\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[27] ),
	.dataf(!\D_src2_reg[27]~45_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[27]~81_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[27]~81 .extended_lut = "off";
defparam \D_src2_reg[27]~81 .lut_mask = 64'hFFFDFFFFFFFFFFFF;
defparam \D_src2_reg[27]~81 .shared_arith = "off";

dffeas \E_src2_reg[27] (
	.clk(clk_clk),
	.d(\D_src2_reg[27]~81_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_src2_reg[27]~q ),
	.prn(vcc));
defparam \E_src2_reg[27] .is_wysiwyg = "true";
defparam \E_src2_reg[27] .power_up = "low";

cyclonev_lcell_comb \E_st_data[27]~5 (
	.dataa(!\E_ctrl_mem16~q ),
	.datab(!\E_src2_reg[11]~q ),
	.datac(!\E_src2_reg[27]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_st_data[27]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_st_data[27]~5 .extended_lut = "off";
defparam \E_st_data[27]~5 .lut_mask = 64'h2727272727272727;
defparam \E_st_data[27]~5 .shared_arith = "off";

dffeas \M_st_data[27] (
	.clk(clk_clk),
	.d(\E_st_data[27]~5_combout ),
	.asdata(\E_src2_reg[3]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_ctrl_mem8~q ),
	.ena(!\A_mem_stall~q ),
	.q(\M_st_data[27]~q ),
	.prn(vcc));
defparam \M_st_data[27] .is_wysiwyg = "true";
defparam \M_st_data[27] .power_up = "low";

dffeas \M_st_data[8] (
	.clk(clk_clk),
	.d(\E_src2_reg[0]~q ),
	.asdata(\E_src2_reg[8]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\E_ctrl_mem8~q ),
	.ena(!\A_mem_stall~q ),
	.q(\M_st_data[8]~q ),
	.prn(vcc));
defparam \M_st_data[8] .is_wysiwyg = "true";
defparam \M_st_data[8] .power_up = "low";

dffeas \M_st_data[9] (
	.clk(clk_clk),
	.d(\E_src2_reg[1]~q ),
	.asdata(\E_src2_reg[9]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\E_ctrl_mem8~q ),
	.ena(!\A_mem_stall~q ),
	.q(\M_st_data[9]~q ),
	.prn(vcc));
defparam \M_st_data[9] .is_wysiwyg = "true";
defparam \M_st_data[9] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[26]~82 (
	.dataa(!\D_src2_reg[26]~53_combout ),
	.datab(!\Equal304~0_combout ),
	.datac(!\D_src2_reg[0]~0_combout ),
	.datad(!\D_src2_reg[0]~1_combout ),
	.datae(!\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[26] ),
	.dataf(!\D_src2_reg[26]~52_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[26]~82_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[26]~82 .extended_lut = "off";
defparam \D_src2_reg[26]~82 .lut_mask = 64'hFFFDFFFFFFFFFFFF;
defparam \D_src2_reg[26]~82 .shared_arith = "off";

dffeas \E_src2_reg[26] (
	.clk(clk_clk),
	.d(\D_src2_reg[26]~82_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_src2_reg[26]~q ),
	.prn(vcc));
defparam \E_src2_reg[26] .is_wysiwyg = "true";
defparam \E_src2_reg[26] .power_up = "low";

cyclonev_lcell_comb \E_st_data[26]~6 (
	.dataa(!\E_ctrl_mem16~q ),
	.datab(!\E_src2_reg[10]~q ),
	.datac(!\E_src2_reg[26]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_st_data[26]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_st_data[26]~6 .extended_lut = "off";
defparam \E_st_data[26]~6 .lut_mask = 64'h2727272727272727;
defparam \E_st_data[26]~6 .shared_arith = "off";

dffeas \M_st_data[26] (
	.clk(clk_clk),
	.d(\E_st_data[26]~6_combout ),
	.asdata(\E_src2_reg[2]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_ctrl_mem8~q ),
	.ena(!\A_mem_stall~q ),
	.q(\M_st_data[26]~q ),
	.prn(vcc));
defparam \M_st_data[26] .is_wysiwyg = "true";
defparam \M_st_data[26] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[20]~83 (
	.dataa(!\D_src2_reg[0]~4_combout ),
	.datab(!\D_src2_reg[0]~5_combout ),
	.datac(!\E_alu_result[20]~combout ),
	.datad(!\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[20] ),
	.datae(!\D_src2_reg[20]~54_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[20]~83_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[20]~83 .extended_lut = "off";
defparam \D_src2_reg[20]~83 .lut_mask = 64'h47FFFFFF47FFFFFF;
defparam \D_src2_reg[20]~83 .shared_arith = "off";

dffeas \E_src2_reg[20] (
	.clk(clk_clk),
	.d(\D_src2_reg[20]~83_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_src2_reg[20]~q ),
	.prn(vcc));
defparam \E_src2_reg[20] .is_wysiwyg = "true";
defparam \E_src2_reg[20] .power_up = "low";

dffeas \M_st_data[20] (
	.clk(clk_clk),
	.d(\E_src2_reg[4]~q ),
	.asdata(\E_src2_reg[20]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_st_data[23]~0_combout ),
	.ena(!\A_mem_stall~q ),
	.q(\M_st_data[20]~q ),
	.prn(vcc));
defparam \M_st_data[20] .is_wysiwyg = "true";
defparam \M_st_data[20] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[19]~84 (
	.dataa(!\D_src2_reg[0]~4_combout ),
	.datab(!\D_src2_reg[0]~5_combout ),
	.datac(!\E_alu_result[19]~combout ),
	.datad(!\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[19] ),
	.datae(!\D_src2_reg[19]~55_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[19]~84_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[19]~84 .extended_lut = "off";
defparam \D_src2_reg[19]~84 .lut_mask = 64'h47FFFFFF47FFFFFF;
defparam \D_src2_reg[19]~84 .shared_arith = "off";

dffeas \E_src2_reg[19] (
	.clk(clk_clk),
	.d(\D_src2_reg[19]~84_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_src2_reg[19]~q ),
	.prn(vcc));
defparam \E_src2_reg[19] .is_wysiwyg = "true";
defparam \E_src2_reg[19] .power_up = "low";

dffeas \M_st_data[19] (
	.clk(clk_clk),
	.d(\E_src2_reg[3]~q ),
	.asdata(\E_src2_reg[19]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_st_data[23]~0_combout ),
	.ena(!\A_mem_stall~q ),
	.q(\M_st_data[19]~q ),
	.prn(vcc));
defparam \M_st_data[19] .is_wysiwyg = "true";
defparam \M_st_data[19] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[17]~85 (
	.dataa(!\D_src2_reg[0]~4_combout ),
	.datab(!\D_src2_reg[0]~5_combout ),
	.datac(!\E_alu_result[17]~combout ),
	.datad(!\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[17] ),
	.datae(!\D_src2_reg[17]~56_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[17]~85_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[17]~85 .extended_lut = "off";
defparam \D_src2_reg[17]~85 .lut_mask = 64'h47FFFFFF47FFFFFF;
defparam \D_src2_reg[17]~85 .shared_arith = "off";

dffeas \E_src2_reg[17] (
	.clk(clk_clk),
	.d(\D_src2_reg[17]~85_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_src2_reg[17]~q ),
	.prn(vcc));
defparam \E_src2_reg[17] .is_wysiwyg = "true";
defparam \E_src2_reg[17] .power_up = "low";

dffeas \M_st_data[17] (
	.clk(clk_clk),
	.d(\E_src2_reg[1]~q ),
	.asdata(\E_src2_reg[17]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_st_data[23]~0_combout ),
	.ena(!\A_mem_stall~q ),
	.q(\M_st_data[17]~q ),
	.prn(vcc));
defparam \M_st_data[17] .is_wysiwyg = "true";
defparam \M_st_data[17] .power_up = "low";

dffeas \E_src2_reg[14] (
	.clk(clk_clk),
	.d(\D_src2_reg[14]~69_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_src2_reg[14]~q ),
	.prn(vcc));
defparam \E_src2_reg[14] .is_wysiwyg = "true";
defparam \E_src2_reg[14] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[30]~86 (
	.dataa(!\D_src2_reg[30]~59_combout ),
	.datab(!\Equal304~0_combout ),
	.datac(!\D_src2_reg[0]~0_combout ),
	.datad(!\D_src2_reg[0]~1_combout ),
	.datae(!\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[30] ),
	.dataf(!\D_src2_reg[30]~57_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[30]~86_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[30]~86 .extended_lut = "off";
defparam \D_src2_reg[30]~86 .lut_mask = 64'hFFFDFFFFFFFFFFFF;
defparam \D_src2_reg[30]~86 .shared_arith = "off";

dffeas \E_src2_reg[30] (
	.clk(clk_clk),
	.d(\D_src2_reg[30]~86_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_src2_reg[30]~q ),
	.prn(vcc));
defparam \E_src2_reg[30] .is_wysiwyg = "true";
defparam \E_src2_reg[30] .power_up = "low";

cyclonev_lcell_comb \E_st_data[30]~7 (
	.dataa(!\E_ctrl_mem16~q ),
	.datab(!\E_src2_reg[14]~q ),
	.datac(!\E_src2_reg[30]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_st_data[30]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_st_data[30]~7 .extended_lut = "off";
defparam \E_st_data[30]~7 .lut_mask = 64'h2727272727272727;
defparam \E_st_data[30]~7 .shared_arith = "off";

dffeas \M_st_data[30] (
	.clk(clk_clk),
	.d(\E_st_data[30]~7_combout ),
	.asdata(\E_src2_reg[6]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_ctrl_mem8~q ),
	.ena(!\A_mem_stall~q ),
	.q(\M_st_data[30]~q ),
	.prn(vcc));
defparam \M_st_data[30] .is_wysiwyg = "true";
defparam \M_st_data[30] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[18]~87 (
	.dataa(!\D_src2_reg[0]~4_combout ),
	.datab(!\D_src2_reg[0]~5_combout ),
	.datac(!\E_alu_result[18]~combout ),
	.datad(!\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[18] ),
	.datae(!\D_src2_reg[18]~60_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[18]~87_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[18]~87 .extended_lut = "off";
defparam \D_src2_reg[18]~87 .lut_mask = 64'h47FFFFFF47FFFFFF;
defparam \D_src2_reg[18]~87 .shared_arith = "off";

dffeas \E_src2_reg[18] (
	.clk(clk_clk),
	.d(\D_src2_reg[18]~87_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_src2_reg[18]~q ),
	.prn(vcc));
defparam \E_src2_reg[18] .is_wysiwyg = "true";
defparam \E_src2_reg[18] .power_up = "low";

dffeas \M_st_data[18] (
	.clk(clk_clk),
	.d(\E_src2_reg[2]~q ),
	.asdata(\E_src2_reg[18]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_st_data[23]~0_combout ),
	.ena(!\A_mem_stall~q ),
	.q(\M_st_data[18]~q ),
	.prn(vcc));
defparam \M_st_data[18] .is_wysiwyg = "true";
defparam \M_st_data[18] .power_up = "low";

dffeas \M_st_data[15] (
	.clk(clk_clk),
	.d(\E_src2_reg[7]~q ),
	.asdata(\E_src2_reg[15]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\E_ctrl_mem8~q ),
	.ena(!\A_mem_stall~q ),
	.q(\M_st_data[15]~q ),
	.prn(vcc));
defparam \M_st_data[15] .is_wysiwyg = "true";
defparam \M_st_data[15] .power_up = "low";

dffeas \M_st_data[12] (
	.clk(clk_clk),
	.d(\E_src2_reg[4]~q ),
	.asdata(\E_src2_reg[12]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\E_ctrl_mem8~q ),
	.ena(!\A_mem_stall~q ),
	.q(\M_st_data[12]~q ),
	.prn(vcc));
defparam \M_st_data[12] .is_wysiwyg = "true";
defparam \M_st_data[12] .power_up = "low";

dffeas \E_src2_reg[13] (
	.clk(clk_clk),
	.d(\D_src2_reg[13]~67_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_src2_reg[13]~q ),
	.prn(vcc));
defparam \E_src2_reg[13] .is_wysiwyg = "true";
defparam \E_src2_reg[13] .power_up = "low";

dffeas \M_st_data[13] (
	.clk(clk_clk),
	.d(\E_src2_reg[5]~q ),
	.asdata(\E_src2_reg[13]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\E_ctrl_mem8~q ),
	.ena(!\A_mem_stall~q ),
	.q(\M_st_data[13]~q ),
	.prn(vcc));
defparam \M_st_data[13] .is_wysiwyg = "true";
defparam \M_st_data[13] .power_up = "low";

dffeas \M_st_data[14] (
	.clk(clk_clk),
	.d(\E_src2_reg[6]~q ),
	.asdata(\E_src2_reg[14]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\E_ctrl_mem8~q ),
	.ena(!\A_mem_stall~q ),
	.q(\M_st_data[14]~q ),
	.prn(vcc));
defparam \M_st_data[14] .is_wysiwyg = "true";
defparam \M_st_data[14] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[29]~88 (
	.dataa(!\D_src2_reg[29]~72_combout ),
	.datab(!\Equal304~0_combout ),
	.datac(!\D_src2_reg[0]~0_combout ),
	.datad(!\D_src2_reg[0]~1_combout ),
	.datae(!\first_nios2_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[29] ),
	.dataf(!\D_src2_reg[29]~70_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[29]~88_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[29]~88 .extended_lut = "off";
defparam \D_src2_reg[29]~88 .lut_mask = 64'hFFFDFFFFFFFFFFFF;
defparam \D_src2_reg[29]~88 .shared_arith = "off";

dffeas \E_src2_reg[29] (
	.clk(clk_clk),
	.d(\D_src2_reg[29]~88_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\A_mem_stall~q ),
	.q(\E_src2_reg[29]~q ),
	.prn(vcc));
defparam \E_src2_reg[29] .is_wysiwyg = "true";
defparam \E_src2_reg[29] .power_up = "low";

cyclonev_lcell_comb \E_st_data[29]~8 (
	.dataa(!\E_ctrl_mem16~q ),
	.datab(!\E_src2_reg[13]~q ),
	.datac(!\E_src2_reg[29]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_st_data[29]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_st_data[29]~8 .extended_lut = "off";
defparam \E_st_data[29]~8 .lut_mask = 64'h2727272727272727;
defparam \E_st_data[29]~8 .shared_arith = "off";

dffeas \M_st_data[29] (
	.clk(clk_clk),
	.d(\E_st_data[29]~8_combout ),
	.asdata(\E_src2_reg[5]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_ctrl_mem8~q ),
	.ena(!\A_mem_stall~q ),
	.q(\M_st_data[29]~q ),
	.prn(vcc));
defparam \M_st_data[29] .is_wysiwyg = "true";
defparam \M_st_data[29] .power_up = "low";

endmodule

module first_nios2_system_first_nios2_system_cpu_cpu_bht_module (
	q_b_1,
	q_b_0,
	F_stall,
	M_bht_wr_en_unfiltered,
	M_bht_wr_data_unfiltered_1,
	M_bht_ptr_unfiltered_0,
	M_bht_ptr_unfiltered_1,
	M_bht_ptr_unfiltered_2,
	M_bht_ptr_unfiltered_3,
	M_bht_ptr_unfiltered_4,
	M_bht_ptr_unfiltered_5,
	M_bht_ptr_unfiltered_6,
	M_bht_ptr_unfiltered_7,
	F_bht_ptr_nxt_0,
	F_bht_ptr_nxt_1,
	F_bht_ptr_nxt_2,
	F_bht_ptr_nxt_3,
	F_bht_ptr_nxt_4,
	F_bht_ptr_nxt_5,
	F_bht_ptr_nxt_6,
	F_bht_ptr_nxt_7,
	M_br_mispredict,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_1;
output 	q_b_0;
input 	F_stall;
input 	M_bht_wr_en_unfiltered;
input 	M_bht_wr_data_unfiltered_1;
input 	M_bht_ptr_unfiltered_0;
input 	M_bht_ptr_unfiltered_1;
input 	M_bht_ptr_unfiltered_2;
input 	M_bht_ptr_unfiltered_3;
input 	M_bht_ptr_unfiltered_4;
input 	M_bht_ptr_unfiltered_5;
input 	M_bht_ptr_unfiltered_6;
input 	M_bht_ptr_unfiltered_7;
input 	F_bht_ptr_nxt_0;
input 	F_bht_ptr_nxt_1;
input 	F_bht_ptr_nxt_2;
input 	F_bht_ptr_nxt_3;
input 	F_bht_ptr_nxt_4;
input 	F_bht_ptr_nxt_5;
input 	F_bht_ptr_nxt_6;
input 	F_bht_ptr_nxt_7;
input 	M_br_mispredict;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



first_nios2_system_altsyncram_1 the_altsyncram(
	.q_b({q_b_unconnected_wire_31,q_b_unconnected_wire_30,q_b_unconnected_wire_29,q_b_unconnected_wire_28,q_b_unconnected_wire_27,q_b_unconnected_wire_26,q_b_unconnected_wire_25,q_b_unconnected_wire_24,q_b_unconnected_wire_23,q_b_unconnected_wire_22,q_b_unconnected_wire_21,
q_b_unconnected_wire_20,q_b_unconnected_wire_19,q_b_unconnected_wire_18,q_b_unconnected_wire_17,q_b_unconnected_wire_16,q_b_unconnected_wire_15,q_b_unconnected_wire_14,q_b_unconnected_wire_13,q_b_unconnected_wire_12,q_b_unconnected_wire_11,q_b_unconnected_wire_10,
q_b_unconnected_wire_9,q_b_unconnected_wire_8,q_b_unconnected_wire_7,q_b_unconnected_wire_6,q_b_unconnected_wire_5,q_b_unconnected_wire_4,q_b_unconnected_wire_3,q_b_unconnected_wire_2,q_b_1,q_b_0}),
	.rden_b(F_stall),
	.wren_a(M_bht_wr_en_unfiltered),
	.data_a({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,M_bht_wr_data_unfiltered_1,M_br_mispredict}),
	.address_a({gnd,gnd,gnd,gnd,gnd,M_bht_ptr_unfiltered_7,M_bht_ptr_unfiltered_6,M_bht_ptr_unfiltered_5,M_bht_ptr_unfiltered_4,M_bht_ptr_unfiltered_3,M_bht_ptr_unfiltered_2,M_bht_ptr_unfiltered_1,M_bht_ptr_unfiltered_0}),
	.address_b({gnd,F_bht_ptr_nxt_7,F_bht_ptr_nxt_6,F_bht_ptr_nxt_5,F_bht_ptr_nxt_4,F_bht_ptr_nxt_3,F_bht_ptr_nxt_2,F_bht_ptr_nxt_1,F_bht_ptr_nxt_0}),
	.clock0(clk_clk));

endmodule

module first_nios2_system_altsyncram_1 (
	q_b,
	rden_b,
	wren_a,
	data_a,
	address_a,
	address_b,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_b;
input 	rden_b;
input 	wren_a;
input 	[31:0] data_a;
input 	[12:0] address_a;
input 	[8:0] address_b;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



first_nios2_system_altsyncram_pdj1 auto_generated(
	.q_b({q_b[1],q_b[0]}),
	.rden_b(rden_b),
	.wren_a(wren_a),
	.data_a({data_a[1],data_a[0]}),
	.address_a({address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.address_b({address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.clock0(clock0));

endmodule

module first_nios2_system_altsyncram_pdj1 (
	q_b,
	rden_b,
	wren_a,
	data_a,
	address_a,
	address_b,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[1:0] q_b;
input 	rden_b;
input 	wren_a;
input 	[1:0] data_a;
input 	[7:0] address_a;
input 	[7:0] address_b;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

cyclonev_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(!rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_bht_module:first_nios2_system_cpu_cpu_bht|altsyncram:the_altsyncram|altsyncram_pdj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "old";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 8;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 255;
defparam ram_block1a1.port_a_logical_ram_depth = 256;
defparam ram_block1a1.port_a_logical_ram_width = 2;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock0";
defparam ram_block1a1.port_b_address_width = 8;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "none";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 255;
defparam ram_block1a1.port_b_logical_ram_depth = 256;
defparam ram_block1a1.port_b_logical_ram_width = 2;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock0";
defparam ram_block1a1.ram_block_type = "auto";

cyclonev_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(!rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_bht_module:first_nios2_system_cpu_cpu_bht|altsyncram:the_altsyncram|altsyncram_pdj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "old";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 8;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 255;
defparam ram_block1a0.port_a_logical_ram_depth = 256;
defparam ram_block1a0.port_a_logical_ram_width = 2;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock0";
defparam ram_block1a0.port_b_address_width = 8;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "none";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 255;
defparam ram_block1a0.port_b_logical_ram_depth = 256;
defparam ram_block1a0.port_b_logical_ram_width = 2;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock0";
defparam ram_block1a0.ram_block_type = "auto";

endmodule

module first_nios2_system_first_nios2_system_cpu_cpu_ic_data_module (
	q_b_26,
	q_b_25,
	q_b_24,
	q_b_23,
	q_b_22,
	q_b_1,
	q_b_0,
	q_b_2,
	q_b_3,
	q_b_4,
	q_b_5,
	q_b_28,
	q_b_31,
	q_b_27,
	q_b_29,
	q_b_30,
	q_b_11,
	q_b_12,
	q_b_13,
	q_b_14,
	q_b_15,
	q_b_16,
	q_b_9,
	q_b_21,
	q_b_6,
	q_b_8,
	q_b_17,
	q_b_18,
	q_b_10,
	q_b_7,
	q_b_20,
	q_b_19,
	ic_fill_line_0,
	ic_fill_line_5,
	ic_fill_line_4,
	ic_fill_line_3,
	ic_fill_line_2,
	ic_fill_line_1,
	F_stall,
	ic_fill_dp_offset_0,
	ic_fill_dp_offset_1,
	ic_fill_dp_offset_2,
	i_readdatavalid_d1,
	i_readdata_d1_26,
	F_ic_data_rd_addr_nxt_0,
	F_ic_data_rd_addr_nxt_1,
	F_ic_data_rd_addr_nxt_2,
	F_ic_tag_rd_addr_nxt_0,
	F_ic_tag_rd_addr_nxt_1,
	F_ic_tag_rd_addr_nxt_2,
	F_ic_tag_rd_addr_nxt_3,
	F_ic_tag_rd_addr_nxt_4,
	F_ic_tag_rd_addr_nxt_5,
	i_readdata_d1_25,
	i_readdata_d1_24,
	i_readdata_d1_23,
	i_readdata_d1_22,
	i_readdata_d1_1,
	i_readdata_d1_0,
	i_readdata_d1_2,
	i_readdata_d1_3,
	i_readdata_d1_4,
	i_readdata_d1_5,
	i_readdata_d1_28,
	i_readdata_d1_31,
	i_readdata_d1_27,
	i_readdata_d1_29,
	i_readdata_d1_30,
	i_readdata_d1_11,
	i_readdata_d1_12,
	i_readdata_d1_13,
	i_readdata_d1_14,
	i_readdata_d1_15,
	i_readdata_d1_16,
	i_readdata_d1_9,
	i_readdata_d1_21,
	i_readdata_d1_6,
	i_readdata_d1_8,
	i_readdata_d1_17,
	i_readdata_d1_18,
	i_readdata_d1_10,
	i_readdata_d1_7,
	i_readdata_d1_20,
	i_readdata_d1_19,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_26;
output 	q_b_25;
output 	q_b_24;
output 	q_b_23;
output 	q_b_22;
output 	q_b_1;
output 	q_b_0;
output 	q_b_2;
output 	q_b_3;
output 	q_b_4;
output 	q_b_5;
output 	q_b_28;
output 	q_b_31;
output 	q_b_27;
output 	q_b_29;
output 	q_b_30;
output 	q_b_11;
output 	q_b_12;
output 	q_b_13;
output 	q_b_14;
output 	q_b_15;
output 	q_b_16;
output 	q_b_9;
output 	q_b_21;
output 	q_b_6;
output 	q_b_8;
output 	q_b_17;
output 	q_b_18;
output 	q_b_10;
output 	q_b_7;
output 	q_b_20;
output 	q_b_19;
input 	ic_fill_line_0;
input 	ic_fill_line_5;
input 	ic_fill_line_4;
input 	ic_fill_line_3;
input 	ic_fill_line_2;
input 	ic_fill_line_1;
input 	F_stall;
input 	ic_fill_dp_offset_0;
input 	ic_fill_dp_offset_1;
input 	ic_fill_dp_offset_2;
input 	i_readdatavalid_d1;
input 	i_readdata_d1_26;
input 	F_ic_data_rd_addr_nxt_0;
input 	F_ic_data_rd_addr_nxt_1;
input 	F_ic_data_rd_addr_nxt_2;
input 	F_ic_tag_rd_addr_nxt_0;
input 	F_ic_tag_rd_addr_nxt_1;
input 	F_ic_tag_rd_addr_nxt_2;
input 	F_ic_tag_rd_addr_nxt_3;
input 	F_ic_tag_rd_addr_nxt_4;
input 	F_ic_tag_rd_addr_nxt_5;
input 	i_readdata_d1_25;
input 	i_readdata_d1_24;
input 	i_readdata_d1_23;
input 	i_readdata_d1_22;
input 	i_readdata_d1_1;
input 	i_readdata_d1_0;
input 	i_readdata_d1_2;
input 	i_readdata_d1_3;
input 	i_readdata_d1_4;
input 	i_readdata_d1_5;
input 	i_readdata_d1_28;
input 	i_readdata_d1_31;
input 	i_readdata_d1_27;
input 	i_readdata_d1_29;
input 	i_readdata_d1_30;
input 	i_readdata_d1_11;
input 	i_readdata_d1_12;
input 	i_readdata_d1_13;
input 	i_readdata_d1_14;
input 	i_readdata_d1_15;
input 	i_readdata_d1_16;
input 	i_readdata_d1_9;
input 	i_readdata_d1_21;
input 	i_readdata_d1_6;
input 	i_readdata_d1_8;
input 	i_readdata_d1_17;
input 	i_readdata_d1_18;
input 	i_readdata_d1_10;
input 	i_readdata_d1_7;
input 	i_readdata_d1_20;
input 	i_readdata_d1_19;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



first_nios2_system_altsyncram_2 the_altsyncram(
	.q_b({q_b_31,q_b_30,q_b_29,q_b_28,q_b_27,q_b_26,q_b_25,q_b_24,q_b_23,q_b_22,q_b_21,q_b_20,q_b_19,q_b_18,q_b_17,q_b_16,q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.address_a({gnd,gnd,gnd,gnd,ic_fill_line_5,ic_fill_line_4,ic_fill_line_3,ic_fill_line_2,ic_fill_line_1,ic_fill_line_0,ic_fill_dp_offset_2,ic_fill_dp_offset_1,ic_fill_dp_offset_0}),
	.rden_b(F_stall),
	.wren_a(i_readdatavalid_d1),
	.data_a({i_readdata_d1_31,i_readdata_d1_30,i_readdata_d1_29,i_readdata_d1_28,i_readdata_d1_27,i_readdata_d1_26,i_readdata_d1_25,i_readdata_d1_24,i_readdata_d1_23,i_readdata_d1_22,i_readdata_d1_21,i_readdata_d1_20,i_readdata_d1_19,i_readdata_d1_18,i_readdata_d1_17,i_readdata_d1_16,
i_readdata_d1_15,i_readdata_d1_14,i_readdata_d1_13,i_readdata_d1_12,i_readdata_d1_11,i_readdata_d1_10,i_readdata_d1_9,i_readdata_d1_8,i_readdata_d1_7,i_readdata_d1_6,i_readdata_d1_5,i_readdata_d1_4,i_readdata_d1_3,i_readdata_d1_2,i_readdata_d1_1,i_readdata_d1_0}),
	.address_b({F_ic_tag_rd_addr_nxt_5,F_ic_tag_rd_addr_nxt_4,F_ic_tag_rd_addr_nxt_3,F_ic_tag_rd_addr_nxt_2,F_ic_tag_rd_addr_nxt_1,F_ic_tag_rd_addr_nxt_0,F_ic_data_rd_addr_nxt_2,F_ic_data_rd_addr_nxt_1,F_ic_data_rd_addr_nxt_0}),
	.clock0(clk_clk));

endmodule

module first_nios2_system_altsyncram_2 (
	q_b,
	address_a,
	rden_b,
	wren_a,
	data_a,
	address_b,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_b;
input 	[12:0] address_a;
input 	rden_b;
input 	wren_a;
input 	[31:0] data_a;
input 	[8:0] address_b;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



first_nios2_system_altsyncram_ekj1 auto_generated(
	.q_b({q_b[31],q_b[30],q_b[29],q_b[28],q_b[27],q_b[26],q_b[25],q_b[24],q_b[23],q_b[22],q_b[21],q_b[20],q_b[19],q_b[18],q_b[17],q_b[16],q_b[15],q_b[14],q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.address_a({address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.rden_b(rden_b),
	.wren_a(wren_a),
	.data_a({data_a[31],data_a[30],data_a[29],data_a[28],data_a[27],data_a[26],data_a[25],data_a[24],data_a[23],data_a[22],data_a[21],data_a[20],data_a[19],data_a[18],data_a[17],data_a[16],data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.address_b({address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.clock0(clock0));

endmodule

module first_nios2_system_altsyncram_ekj1 (
	q_b,
	address_a,
	rden_b,
	wren_a,
	data_a,
	address_b,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_b;
input 	[8:0] address_a;
input 	rden_b;
input 	wren_a;
input 	[31:0] data_a;
input 	[8:0] address_b;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a26_PORTBDATAOUT_bus;
wire [143:0] ram_block1a25_PORTBDATAOUT_bus;
wire [143:0] ram_block1a24_PORTBDATAOUT_bus;
wire [143:0] ram_block1a23_PORTBDATAOUT_bus;
wire [143:0] ram_block1a22_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a28_PORTBDATAOUT_bus;
wire [143:0] ram_block1a31_PORTBDATAOUT_bus;
wire [143:0] ram_block1a27_PORTBDATAOUT_bus;
wire [143:0] ram_block1a29_PORTBDATAOUT_bus;
wire [143:0] ram_block1a30_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a21_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a20_PORTBDATAOUT_bus;
wire [143:0] ram_block1a19_PORTBDATAOUT_bus;

assign q_b[26] = ram_block1a26_PORTBDATAOUT_bus[0];

assign q_b[25] = ram_block1a25_PORTBDATAOUT_bus[0];

assign q_b[24] = ram_block1a24_PORTBDATAOUT_bus[0];

assign q_b[23] = ram_block1a23_PORTBDATAOUT_bus[0];

assign q_b[22] = ram_block1a22_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[28] = ram_block1a28_PORTBDATAOUT_bus[0];

assign q_b[31] = ram_block1a31_PORTBDATAOUT_bus[0];

assign q_b[27] = ram_block1a27_PORTBDATAOUT_bus[0];

assign q_b[29] = ram_block1a29_PORTBDATAOUT_bus[0];

assign q_b[30] = ram_block1a30_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[16] = ram_block1a16_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[21] = ram_block1a21_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[17] = ram_block1a17_PORTBDATAOUT_bus[0];

assign q_b[18] = ram_block1a18_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[20] = ram_block1a20_PORTBDATAOUT_bus[0];

assign q_b[19] = ram_block1a19_PORTBDATAOUT_bus[0];

cyclonev_ram_block ram_block1a26(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[26]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a26_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a26.clk0_core_clock_enable = "ena0";
defparam ram_block1a26.clk1_core_clock_enable = "ena1";
defparam ram_block1a26.data_interleave_offset_in_bits = 1;
defparam ram_block1a26.data_interleave_width_in_bits = 1;
defparam ram_block1a26.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_ic_data_module:first_nios2_system_cpu_cpu_ic_data|altsyncram:the_altsyncram|altsyncram_ekj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a26.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a26.operation_mode = "dual_port";
defparam ram_block1a26.port_a_address_clear = "none";
defparam ram_block1a26.port_a_address_width = 9;
defparam ram_block1a26.port_a_data_out_clear = "none";
defparam ram_block1a26.port_a_data_out_clock = "none";
defparam ram_block1a26.port_a_data_width = 1;
defparam ram_block1a26.port_a_first_address = 0;
defparam ram_block1a26.port_a_first_bit_number = 26;
defparam ram_block1a26.port_a_last_address = 511;
defparam ram_block1a26.port_a_logical_ram_depth = 512;
defparam ram_block1a26.port_a_logical_ram_width = 32;
defparam ram_block1a26.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a26.port_b_address_clear = "none";
defparam ram_block1a26.port_b_address_clock = "clock1";
defparam ram_block1a26.port_b_address_width = 9;
defparam ram_block1a26.port_b_data_out_clear = "none";
defparam ram_block1a26.port_b_data_out_clock = "none";
defparam ram_block1a26.port_b_data_width = 1;
defparam ram_block1a26.port_b_first_address = 0;
defparam ram_block1a26.port_b_first_bit_number = 26;
defparam ram_block1a26.port_b_last_address = 511;
defparam ram_block1a26.port_b_logical_ram_depth = 512;
defparam ram_block1a26.port_b_logical_ram_width = 32;
defparam ram_block1a26.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a26.port_b_read_enable_clock = "clock1";
defparam ram_block1a26.ram_block_type = "auto";

cyclonev_ram_block ram_block1a25(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[25]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a25_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a25.clk0_core_clock_enable = "ena0";
defparam ram_block1a25.clk1_core_clock_enable = "ena1";
defparam ram_block1a25.data_interleave_offset_in_bits = 1;
defparam ram_block1a25.data_interleave_width_in_bits = 1;
defparam ram_block1a25.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_ic_data_module:first_nios2_system_cpu_cpu_ic_data|altsyncram:the_altsyncram|altsyncram_ekj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a25.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a25.operation_mode = "dual_port";
defparam ram_block1a25.port_a_address_clear = "none";
defparam ram_block1a25.port_a_address_width = 9;
defparam ram_block1a25.port_a_data_out_clear = "none";
defparam ram_block1a25.port_a_data_out_clock = "none";
defparam ram_block1a25.port_a_data_width = 1;
defparam ram_block1a25.port_a_first_address = 0;
defparam ram_block1a25.port_a_first_bit_number = 25;
defparam ram_block1a25.port_a_last_address = 511;
defparam ram_block1a25.port_a_logical_ram_depth = 512;
defparam ram_block1a25.port_a_logical_ram_width = 32;
defparam ram_block1a25.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a25.port_b_address_clear = "none";
defparam ram_block1a25.port_b_address_clock = "clock1";
defparam ram_block1a25.port_b_address_width = 9;
defparam ram_block1a25.port_b_data_out_clear = "none";
defparam ram_block1a25.port_b_data_out_clock = "none";
defparam ram_block1a25.port_b_data_width = 1;
defparam ram_block1a25.port_b_first_address = 0;
defparam ram_block1a25.port_b_first_bit_number = 25;
defparam ram_block1a25.port_b_last_address = 511;
defparam ram_block1a25.port_b_logical_ram_depth = 512;
defparam ram_block1a25.port_b_logical_ram_width = 32;
defparam ram_block1a25.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a25.port_b_read_enable_clock = "clock1";
defparam ram_block1a25.ram_block_type = "auto";

cyclonev_ram_block ram_block1a24(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[24]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a24_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a24.clk0_core_clock_enable = "ena0";
defparam ram_block1a24.clk1_core_clock_enable = "ena1";
defparam ram_block1a24.data_interleave_offset_in_bits = 1;
defparam ram_block1a24.data_interleave_width_in_bits = 1;
defparam ram_block1a24.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_ic_data_module:first_nios2_system_cpu_cpu_ic_data|altsyncram:the_altsyncram|altsyncram_ekj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a24.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a24.operation_mode = "dual_port";
defparam ram_block1a24.port_a_address_clear = "none";
defparam ram_block1a24.port_a_address_width = 9;
defparam ram_block1a24.port_a_data_out_clear = "none";
defparam ram_block1a24.port_a_data_out_clock = "none";
defparam ram_block1a24.port_a_data_width = 1;
defparam ram_block1a24.port_a_first_address = 0;
defparam ram_block1a24.port_a_first_bit_number = 24;
defparam ram_block1a24.port_a_last_address = 511;
defparam ram_block1a24.port_a_logical_ram_depth = 512;
defparam ram_block1a24.port_a_logical_ram_width = 32;
defparam ram_block1a24.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a24.port_b_address_clear = "none";
defparam ram_block1a24.port_b_address_clock = "clock1";
defparam ram_block1a24.port_b_address_width = 9;
defparam ram_block1a24.port_b_data_out_clear = "none";
defparam ram_block1a24.port_b_data_out_clock = "none";
defparam ram_block1a24.port_b_data_width = 1;
defparam ram_block1a24.port_b_first_address = 0;
defparam ram_block1a24.port_b_first_bit_number = 24;
defparam ram_block1a24.port_b_last_address = 511;
defparam ram_block1a24.port_b_logical_ram_depth = 512;
defparam ram_block1a24.port_b_logical_ram_width = 32;
defparam ram_block1a24.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a24.port_b_read_enable_clock = "clock1";
defparam ram_block1a24.ram_block_type = "auto";

cyclonev_ram_block ram_block1a23(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[23]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a23_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a23.clk0_core_clock_enable = "ena0";
defparam ram_block1a23.clk1_core_clock_enable = "ena1";
defparam ram_block1a23.data_interleave_offset_in_bits = 1;
defparam ram_block1a23.data_interleave_width_in_bits = 1;
defparam ram_block1a23.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_ic_data_module:first_nios2_system_cpu_cpu_ic_data|altsyncram:the_altsyncram|altsyncram_ekj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a23.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a23.operation_mode = "dual_port";
defparam ram_block1a23.port_a_address_clear = "none";
defparam ram_block1a23.port_a_address_width = 9;
defparam ram_block1a23.port_a_data_out_clear = "none";
defparam ram_block1a23.port_a_data_out_clock = "none";
defparam ram_block1a23.port_a_data_width = 1;
defparam ram_block1a23.port_a_first_address = 0;
defparam ram_block1a23.port_a_first_bit_number = 23;
defparam ram_block1a23.port_a_last_address = 511;
defparam ram_block1a23.port_a_logical_ram_depth = 512;
defparam ram_block1a23.port_a_logical_ram_width = 32;
defparam ram_block1a23.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a23.port_b_address_clear = "none";
defparam ram_block1a23.port_b_address_clock = "clock1";
defparam ram_block1a23.port_b_address_width = 9;
defparam ram_block1a23.port_b_data_out_clear = "none";
defparam ram_block1a23.port_b_data_out_clock = "none";
defparam ram_block1a23.port_b_data_width = 1;
defparam ram_block1a23.port_b_first_address = 0;
defparam ram_block1a23.port_b_first_bit_number = 23;
defparam ram_block1a23.port_b_last_address = 511;
defparam ram_block1a23.port_b_logical_ram_depth = 512;
defparam ram_block1a23.port_b_logical_ram_width = 32;
defparam ram_block1a23.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a23.port_b_read_enable_clock = "clock1";
defparam ram_block1a23.ram_block_type = "auto";

cyclonev_ram_block ram_block1a22(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[22]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a22_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a22.clk0_core_clock_enable = "ena0";
defparam ram_block1a22.clk1_core_clock_enable = "ena1";
defparam ram_block1a22.data_interleave_offset_in_bits = 1;
defparam ram_block1a22.data_interleave_width_in_bits = 1;
defparam ram_block1a22.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_ic_data_module:first_nios2_system_cpu_cpu_ic_data|altsyncram:the_altsyncram|altsyncram_ekj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a22.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a22.operation_mode = "dual_port";
defparam ram_block1a22.port_a_address_clear = "none";
defparam ram_block1a22.port_a_address_width = 9;
defparam ram_block1a22.port_a_data_out_clear = "none";
defparam ram_block1a22.port_a_data_out_clock = "none";
defparam ram_block1a22.port_a_data_width = 1;
defparam ram_block1a22.port_a_first_address = 0;
defparam ram_block1a22.port_a_first_bit_number = 22;
defparam ram_block1a22.port_a_last_address = 511;
defparam ram_block1a22.port_a_logical_ram_depth = 512;
defparam ram_block1a22.port_a_logical_ram_width = 32;
defparam ram_block1a22.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a22.port_b_address_clear = "none";
defparam ram_block1a22.port_b_address_clock = "clock1";
defparam ram_block1a22.port_b_address_width = 9;
defparam ram_block1a22.port_b_data_out_clear = "none";
defparam ram_block1a22.port_b_data_out_clock = "none";
defparam ram_block1a22.port_b_data_width = 1;
defparam ram_block1a22.port_b_first_address = 0;
defparam ram_block1a22.port_b_first_bit_number = 22;
defparam ram_block1a22.port_b_last_address = 511;
defparam ram_block1a22.port_b_logical_ram_depth = 512;
defparam ram_block1a22.port_b_logical_ram_width = 32;
defparam ram_block1a22.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a22.port_b_read_enable_clock = "clock1";
defparam ram_block1a22.ram_block_type = "auto";

cyclonev_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk1_core_clock_enable = "ena1";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_ic_data_module:first_nios2_system_cpu_cpu_ic_data|altsyncram:the_altsyncram|altsyncram_ekj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 9;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 511;
defparam ram_block1a1.port_a_logical_ram_depth = 512;
defparam ram_block1a1.port_a_logical_ram_width = 32;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock1";
defparam ram_block1a1.port_b_address_width = 9;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "none";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 511;
defparam ram_block1a1.port_b_logical_ram_depth = 512;
defparam ram_block1a1.port_b_logical_ram_width = 32;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock1";
defparam ram_block1a1.ram_block_type = "auto";

cyclonev_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk1_core_clock_enable = "ena1";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_ic_data_module:first_nios2_system_cpu_cpu_ic_data|altsyncram:the_altsyncram|altsyncram_ekj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 9;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 511;
defparam ram_block1a0.port_a_logical_ram_depth = 512;
defparam ram_block1a0.port_a_logical_ram_width = 32;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock1";
defparam ram_block1a0.port_b_address_width = 9;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "none";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 511;
defparam ram_block1a0.port_b_logical_ram_depth = 512;
defparam ram_block1a0.port_b_logical_ram_width = 32;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock1";
defparam ram_block1a0.ram_block_type = "auto";

cyclonev_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk1_core_clock_enable = "ena1";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_ic_data_module:first_nios2_system_cpu_cpu_ic_data|altsyncram:the_altsyncram|altsyncram_ekj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 9;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 511;
defparam ram_block1a2.port_a_logical_ram_depth = 512;
defparam ram_block1a2.port_a_logical_ram_width = 32;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock1";
defparam ram_block1a2.port_b_address_width = 9;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "none";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 511;
defparam ram_block1a2.port_b_logical_ram_depth = 512;
defparam ram_block1a2.port_b_logical_ram_width = 32;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock1";
defparam ram_block1a2.ram_block_type = "auto";

cyclonev_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk1_core_clock_enable = "ena1";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_ic_data_module:first_nios2_system_cpu_cpu_ic_data|altsyncram:the_altsyncram|altsyncram_ekj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 9;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 511;
defparam ram_block1a3.port_a_logical_ram_depth = 512;
defparam ram_block1a3.port_a_logical_ram_width = 32;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock1";
defparam ram_block1a3.port_b_address_width = 9;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "none";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 511;
defparam ram_block1a3.port_b_logical_ram_depth = 512;
defparam ram_block1a3.port_b_logical_ram_width = 32;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock1";
defparam ram_block1a3.ram_block_type = "auto";

cyclonev_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk1_core_clock_enable = "ena1";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_ic_data_module:first_nios2_system_cpu_cpu_ic_data|altsyncram:the_altsyncram|altsyncram_ekj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 9;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 511;
defparam ram_block1a4.port_a_logical_ram_depth = 512;
defparam ram_block1a4.port_a_logical_ram_width = 32;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock1";
defparam ram_block1a4.port_b_address_width = 9;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "none";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 511;
defparam ram_block1a4.port_b_logical_ram_depth = 512;
defparam ram_block1a4.port_b_logical_ram_width = 32;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock1";
defparam ram_block1a4.ram_block_type = "auto";

cyclonev_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk1_core_clock_enable = "ena1";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_ic_data_module:first_nios2_system_cpu_cpu_ic_data|altsyncram:the_altsyncram|altsyncram_ekj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 9;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 511;
defparam ram_block1a5.port_a_logical_ram_depth = 512;
defparam ram_block1a5.port_a_logical_ram_width = 32;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 9;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "none";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 511;
defparam ram_block1a5.port_b_logical_ram_depth = 512;
defparam ram_block1a5.port_b_logical_ram_width = 32;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";

cyclonev_ram_block ram_block1a28(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[28]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a28_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a28.clk0_core_clock_enable = "ena0";
defparam ram_block1a28.clk1_core_clock_enable = "ena1";
defparam ram_block1a28.data_interleave_offset_in_bits = 1;
defparam ram_block1a28.data_interleave_width_in_bits = 1;
defparam ram_block1a28.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_ic_data_module:first_nios2_system_cpu_cpu_ic_data|altsyncram:the_altsyncram|altsyncram_ekj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a28.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a28.operation_mode = "dual_port";
defparam ram_block1a28.port_a_address_clear = "none";
defparam ram_block1a28.port_a_address_width = 9;
defparam ram_block1a28.port_a_data_out_clear = "none";
defparam ram_block1a28.port_a_data_out_clock = "none";
defparam ram_block1a28.port_a_data_width = 1;
defparam ram_block1a28.port_a_first_address = 0;
defparam ram_block1a28.port_a_first_bit_number = 28;
defparam ram_block1a28.port_a_last_address = 511;
defparam ram_block1a28.port_a_logical_ram_depth = 512;
defparam ram_block1a28.port_a_logical_ram_width = 32;
defparam ram_block1a28.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a28.port_b_address_clear = "none";
defparam ram_block1a28.port_b_address_clock = "clock1";
defparam ram_block1a28.port_b_address_width = 9;
defparam ram_block1a28.port_b_data_out_clear = "none";
defparam ram_block1a28.port_b_data_out_clock = "none";
defparam ram_block1a28.port_b_data_width = 1;
defparam ram_block1a28.port_b_first_address = 0;
defparam ram_block1a28.port_b_first_bit_number = 28;
defparam ram_block1a28.port_b_last_address = 511;
defparam ram_block1a28.port_b_logical_ram_depth = 512;
defparam ram_block1a28.port_b_logical_ram_width = 32;
defparam ram_block1a28.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a28.port_b_read_enable_clock = "clock1";
defparam ram_block1a28.ram_block_type = "auto";

cyclonev_ram_block ram_block1a31(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a31_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a31.clk0_core_clock_enable = "ena0";
defparam ram_block1a31.clk1_core_clock_enable = "ena1";
defparam ram_block1a31.data_interleave_offset_in_bits = 1;
defparam ram_block1a31.data_interleave_width_in_bits = 1;
defparam ram_block1a31.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_ic_data_module:first_nios2_system_cpu_cpu_ic_data|altsyncram:the_altsyncram|altsyncram_ekj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a31.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a31.operation_mode = "dual_port";
defparam ram_block1a31.port_a_address_clear = "none";
defparam ram_block1a31.port_a_address_width = 9;
defparam ram_block1a31.port_a_data_out_clear = "none";
defparam ram_block1a31.port_a_data_out_clock = "none";
defparam ram_block1a31.port_a_data_width = 1;
defparam ram_block1a31.port_a_first_address = 0;
defparam ram_block1a31.port_a_first_bit_number = 31;
defparam ram_block1a31.port_a_last_address = 511;
defparam ram_block1a31.port_a_logical_ram_depth = 512;
defparam ram_block1a31.port_a_logical_ram_width = 32;
defparam ram_block1a31.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a31.port_b_address_clear = "none";
defparam ram_block1a31.port_b_address_clock = "clock1";
defparam ram_block1a31.port_b_address_width = 9;
defparam ram_block1a31.port_b_data_out_clear = "none";
defparam ram_block1a31.port_b_data_out_clock = "none";
defparam ram_block1a31.port_b_data_width = 1;
defparam ram_block1a31.port_b_first_address = 0;
defparam ram_block1a31.port_b_first_bit_number = 31;
defparam ram_block1a31.port_b_last_address = 511;
defparam ram_block1a31.port_b_logical_ram_depth = 512;
defparam ram_block1a31.port_b_logical_ram_width = 32;
defparam ram_block1a31.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a31.port_b_read_enable_clock = "clock1";
defparam ram_block1a31.ram_block_type = "auto";

cyclonev_ram_block ram_block1a27(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[27]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a27_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a27.clk0_core_clock_enable = "ena0";
defparam ram_block1a27.clk1_core_clock_enable = "ena1";
defparam ram_block1a27.data_interleave_offset_in_bits = 1;
defparam ram_block1a27.data_interleave_width_in_bits = 1;
defparam ram_block1a27.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_ic_data_module:first_nios2_system_cpu_cpu_ic_data|altsyncram:the_altsyncram|altsyncram_ekj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a27.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a27.operation_mode = "dual_port";
defparam ram_block1a27.port_a_address_clear = "none";
defparam ram_block1a27.port_a_address_width = 9;
defparam ram_block1a27.port_a_data_out_clear = "none";
defparam ram_block1a27.port_a_data_out_clock = "none";
defparam ram_block1a27.port_a_data_width = 1;
defparam ram_block1a27.port_a_first_address = 0;
defparam ram_block1a27.port_a_first_bit_number = 27;
defparam ram_block1a27.port_a_last_address = 511;
defparam ram_block1a27.port_a_logical_ram_depth = 512;
defparam ram_block1a27.port_a_logical_ram_width = 32;
defparam ram_block1a27.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a27.port_b_address_clear = "none";
defparam ram_block1a27.port_b_address_clock = "clock1";
defparam ram_block1a27.port_b_address_width = 9;
defparam ram_block1a27.port_b_data_out_clear = "none";
defparam ram_block1a27.port_b_data_out_clock = "none";
defparam ram_block1a27.port_b_data_width = 1;
defparam ram_block1a27.port_b_first_address = 0;
defparam ram_block1a27.port_b_first_bit_number = 27;
defparam ram_block1a27.port_b_last_address = 511;
defparam ram_block1a27.port_b_logical_ram_depth = 512;
defparam ram_block1a27.port_b_logical_ram_width = 32;
defparam ram_block1a27.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a27.port_b_read_enable_clock = "clock1";
defparam ram_block1a27.ram_block_type = "auto";

cyclonev_ram_block ram_block1a29(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[29]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a29_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a29.clk0_core_clock_enable = "ena0";
defparam ram_block1a29.clk1_core_clock_enable = "ena1";
defparam ram_block1a29.data_interleave_offset_in_bits = 1;
defparam ram_block1a29.data_interleave_width_in_bits = 1;
defparam ram_block1a29.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_ic_data_module:first_nios2_system_cpu_cpu_ic_data|altsyncram:the_altsyncram|altsyncram_ekj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a29.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a29.operation_mode = "dual_port";
defparam ram_block1a29.port_a_address_clear = "none";
defparam ram_block1a29.port_a_address_width = 9;
defparam ram_block1a29.port_a_data_out_clear = "none";
defparam ram_block1a29.port_a_data_out_clock = "none";
defparam ram_block1a29.port_a_data_width = 1;
defparam ram_block1a29.port_a_first_address = 0;
defparam ram_block1a29.port_a_first_bit_number = 29;
defparam ram_block1a29.port_a_last_address = 511;
defparam ram_block1a29.port_a_logical_ram_depth = 512;
defparam ram_block1a29.port_a_logical_ram_width = 32;
defparam ram_block1a29.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a29.port_b_address_clear = "none";
defparam ram_block1a29.port_b_address_clock = "clock1";
defparam ram_block1a29.port_b_address_width = 9;
defparam ram_block1a29.port_b_data_out_clear = "none";
defparam ram_block1a29.port_b_data_out_clock = "none";
defparam ram_block1a29.port_b_data_width = 1;
defparam ram_block1a29.port_b_first_address = 0;
defparam ram_block1a29.port_b_first_bit_number = 29;
defparam ram_block1a29.port_b_last_address = 511;
defparam ram_block1a29.port_b_logical_ram_depth = 512;
defparam ram_block1a29.port_b_logical_ram_width = 32;
defparam ram_block1a29.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a29.port_b_read_enable_clock = "clock1";
defparam ram_block1a29.ram_block_type = "auto";

cyclonev_ram_block ram_block1a30(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[30]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a30_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a30.clk0_core_clock_enable = "ena0";
defparam ram_block1a30.clk1_core_clock_enable = "ena1";
defparam ram_block1a30.data_interleave_offset_in_bits = 1;
defparam ram_block1a30.data_interleave_width_in_bits = 1;
defparam ram_block1a30.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_ic_data_module:first_nios2_system_cpu_cpu_ic_data|altsyncram:the_altsyncram|altsyncram_ekj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a30.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a30.operation_mode = "dual_port";
defparam ram_block1a30.port_a_address_clear = "none";
defparam ram_block1a30.port_a_address_width = 9;
defparam ram_block1a30.port_a_data_out_clear = "none";
defparam ram_block1a30.port_a_data_out_clock = "none";
defparam ram_block1a30.port_a_data_width = 1;
defparam ram_block1a30.port_a_first_address = 0;
defparam ram_block1a30.port_a_first_bit_number = 30;
defparam ram_block1a30.port_a_last_address = 511;
defparam ram_block1a30.port_a_logical_ram_depth = 512;
defparam ram_block1a30.port_a_logical_ram_width = 32;
defparam ram_block1a30.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a30.port_b_address_clear = "none";
defparam ram_block1a30.port_b_address_clock = "clock1";
defparam ram_block1a30.port_b_address_width = 9;
defparam ram_block1a30.port_b_data_out_clear = "none";
defparam ram_block1a30.port_b_data_out_clock = "none";
defparam ram_block1a30.port_b_data_width = 1;
defparam ram_block1a30.port_b_first_address = 0;
defparam ram_block1a30.port_b_first_bit_number = 30;
defparam ram_block1a30.port_b_last_address = 511;
defparam ram_block1a30.port_b_logical_ram_depth = 512;
defparam ram_block1a30.port_b_logical_ram_width = 32;
defparam ram_block1a30.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a30.port_b_read_enable_clock = "clock1";
defparam ram_block1a30.ram_block_type = "auto";

cyclonev_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.clk1_core_clock_enable = "ena1";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_ic_data_module:first_nios2_system_cpu_cpu_ic_data|altsyncram:the_altsyncram|altsyncram_ekj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 9;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 511;
defparam ram_block1a11.port_a_logical_ram_depth = 512;
defparam ram_block1a11.port_a_logical_ram_width = 32;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock1";
defparam ram_block1a11.port_b_address_width = 9;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "none";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 511;
defparam ram_block1a11.port_b_logical_ram_depth = 512;
defparam ram_block1a11.port_b_logical_ram_width = 32;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock1";
defparam ram_block1a11.ram_block_type = "auto";

cyclonev_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.clk1_core_clock_enable = "ena1";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_ic_data_module:first_nios2_system_cpu_cpu_ic_data|altsyncram:the_altsyncram|altsyncram_ekj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 9;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 511;
defparam ram_block1a12.port_a_logical_ram_depth = 512;
defparam ram_block1a12.port_a_logical_ram_width = 32;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock1";
defparam ram_block1a12.port_b_address_width = 9;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "none";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 511;
defparam ram_block1a12.port_b_logical_ram_depth = 512;
defparam ram_block1a12.port_b_logical_ram_width = 32;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock1";
defparam ram_block1a12.ram_block_type = "auto";

cyclonev_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.clk1_core_clock_enable = "ena1";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_ic_data_module:first_nios2_system_cpu_cpu_ic_data|altsyncram:the_altsyncram|altsyncram_ekj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 9;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 511;
defparam ram_block1a13.port_a_logical_ram_depth = 512;
defparam ram_block1a13.port_a_logical_ram_width = 32;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock1";
defparam ram_block1a13.port_b_address_width = 9;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "none";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 511;
defparam ram_block1a13.port_b_logical_ram_depth = 512;
defparam ram_block1a13.port_b_logical_ram_width = 32;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock1";
defparam ram_block1a13.ram_block_type = "auto";

cyclonev_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.clk1_core_clock_enable = "ena1";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_ic_data_module:first_nios2_system_cpu_cpu_ic_data|altsyncram:the_altsyncram|altsyncram_ekj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 9;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 511;
defparam ram_block1a14.port_a_logical_ram_depth = 512;
defparam ram_block1a14.port_a_logical_ram_width = 32;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock1";
defparam ram_block1a14.port_b_address_width = 9;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "none";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 511;
defparam ram_block1a14.port_b_logical_ram_depth = 512;
defparam ram_block1a14.port_b_logical_ram_width = 32;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock1";
defparam ram_block1a14.ram_block_type = "auto";

cyclonev_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.clk1_core_clock_enable = "ena1";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_ic_data_module:first_nios2_system_cpu_cpu_ic_data|altsyncram:the_altsyncram|altsyncram_ekj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 9;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 511;
defparam ram_block1a15.port_a_logical_ram_depth = 512;
defparam ram_block1a15.port_a_logical_ram_width = 32;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock1";
defparam ram_block1a15.port_b_address_width = 9;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "none";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 511;
defparam ram_block1a15.port_b_logical_ram_depth = 512;
defparam ram_block1a15.port_b_logical_ram_width = 32;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock1";
defparam ram_block1a15.ram_block_type = "auto";

cyclonev_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a16.clk0_core_clock_enable = "ena0";
defparam ram_block1a16.clk1_core_clock_enable = "ena1";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_ic_data_module:first_nios2_system_cpu_cpu_ic_data|altsyncram:the_altsyncram|altsyncram_ekj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a16.operation_mode = "dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 9;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 511;
defparam ram_block1a16.port_a_logical_ram_depth = 512;
defparam ram_block1a16.port_a_logical_ram_width = 32;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a16.port_b_address_clear = "none";
defparam ram_block1a16.port_b_address_clock = "clock1";
defparam ram_block1a16.port_b_address_width = 9;
defparam ram_block1a16.port_b_data_out_clear = "none";
defparam ram_block1a16.port_b_data_out_clock = "none";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 511;
defparam ram_block1a16.port_b_logical_ram_depth = 512;
defparam ram_block1a16.port_b_logical_ram_width = 32;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock1";
defparam ram_block1a16.ram_block_type = "auto";

cyclonev_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk1_core_clock_enable = "ena1";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_ic_data_module:first_nios2_system_cpu_cpu_ic_data|altsyncram:the_altsyncram|altsyncram_ekj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 9;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 511;
defparam ram_block1a9.port_a_logical_ram_depth = 512;
defparam ram_block1a9.port_a_logical_ram_width = 32;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock1";
defparam ram_block1a9.port_b_address_width = 9;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "none";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 511;
defparam ram_block1a9.port_b_logical_ram_depth = 512;
defparam ram_block1a9.port_b_logical_ram_width = 32;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock1";
defparam ram_block1a9.ram_block_type = "auto";

cyclonev_ram_block ram_block1a21(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a21_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a21.clk0_core_clock_enable = "ena0";
defparam ram_block1a21.clk1_core_clock_enable = "ena1";
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_ic_data_module:first_nios2_system_cpu_cpu_ic_data|altsyncram:the_altsyncram|altsyncram_ekj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a21.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a21.operation_mode = "dual_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 9;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 511;
defparam ram_block1a21.port_a_logical_ram_depth = 512;
defparam ram_block1a21.port_a_logical_ram_width = 32;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a21.port_b_address_clear = "none";
defparam ram_block1a21.port_b_address_clock = "clock1";
defparam ram_block1a21.port_b_address_width = 9;
defparam ram_block1a21.port_b_data_out_clear = "none";
defparam ram_block1a21.port_b_data_out_clock = "none";
defparam ram_block1a21.port_b_data_width = 1;
defparam ram_block1a21.port_b_first_address = 0;
defparam ram_block1a21.port_b_first_bit_number = 21;
defparam ram_block1a21.port_b_last_address = 511;
defparam ram_block1a21.port_b_logical_ram_depth = 512;
defparam ram_block1a21.port_b_logical_ram_width = 32;
defparam ram_block1a21.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a21.port_b_read_enable_clock = "clock1";
defparam ram_block1a21.ram_block_type = "auto";

cyclonev_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk1_core_clock_enable = "ena1";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_ic_data_module:first_nios2_system_cpu_cpu_ic_data|altsyncram:the_altsyncram|altsyncram_ekj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 9;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 511;
defparam ram_block1a6.port_a_logical_ram_depth = 512;
defparam ram_block1a6.port_a_logical_ram_width = 32;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 9;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "none";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 511;
defparam ram_block1a6.port_b_logical_ram_depth = 512;
defparam ram_block1a6.port_b_logical_ram_width = 32;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";

cyclonev_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk1_core_clock_enable = "ena1";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_ic_data_module:first_nios2_system_cpu_cpu_ic_data|altsyncram:the_altsyncram|altsyncram_ekj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 9;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 511;
defparam ram_block1a8.port_a_logical_ram_depth = 512;
defparam ram_block1a8.port_a_logical_ram_width = 32;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock1";
defparam ram_block1a8.port_b_address_width = 9;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "none";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 511;
defparam ram_block1a8.port_b_logical_ram_depth = 512;
defparam ram_block1a8.port_b_logical_ram_width = 32;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock1";
defparam ram_block1a8.ram_block_type = "auto";

cyclonev_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a17.clk0_core_clock_enable = "ena0";
defparam ram_block1a17.clk1_core_clock_enable = "ena1";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_ic_data_module:first_nios2_system_cpu_cpu_ic_data|altsyncram:the_altsyncram|altsyncram_ekj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a17.operation_mode = "dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 9;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 511;
defparam ram_block1a17.port_a_logical_ram_depth = 512;
defparam ram_block1a17.port_a_logical_ram_width = 32;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a17.port_b_address_clear = "none";
defparam ram_block1a17.port_b_address_clock = "clock1";
defparam ram_block1a17.port_b_address_width = 9;
defparam ram_block1a17.port_b_data_out_clear = "none";
defparam ram_block1a17.port_b_data_out_clock = "none";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 511;
defparam ram_block1a17.port_b_logical_ram_depth = 512;
defparam ram_block1a17.port_b_logical_ram_width = 32;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock1";
defparam ram_block1a17.ram_block_type = "auto";

cyclonev_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a18.clk0_core_clock_enable = "ena0";
defparam ram_block1a18.clk1_core_clock_enable = "ena1";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_ic_data_module:first_nios2_system_cpu_cpu_ic_data|altsyncram:the_altsyncram|altsyncram_ekj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a18.operation_mode = "dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 9;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 511;
defparam ram_block1a18.port_a_logical_ram_depth = 512;
defparam ram_block1a18.port_a_logical_ram_width = 32;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a18.port_b_address_clear = "none";
defparam ram_block1a18.port_b_address_clock = "clock1";
defparam ram_block1a18.port_b_address_width = 9;
defparam ram_block1a18.port_b_data_out_clear = "none";
defparam ram_block1a18.port_b_data_out_clock = "none";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 511;
defparam ram_block1a18.port_b_logical_ram_depth = 512;
defparam ram_block1a18.port_b_logical_ram_width = 32;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock1";
defparam ram_block1a18.ram_block_type = "auto";

cyclonev_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.clk1_core_clock_enable = "ena1";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_ic_data_module:first_nios2_system_cpu_cpu_ic_data|altsyncram:the_altsyncram|altsyncram_ekj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 9;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 511;
defparam ram_block1a10.port_a_logical_ram_depth = 512;
defparam ram_block1a10.port_a_logical_ram_width = 32;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock1";
defparam ram_block1a10.port_b_address_width = 9;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "none";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 511;
defparam ram_block1a10.port_b_logical_ram_depth = 512;
defparam ram_block1a10.port_b_logical_ram_width = 32;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock1";
defparam ram_block1a10.ram_block_type = "auto";

cyclonev_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk1_core_clock_enable = "ena1";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_ic_data_module:first_nios2_system_cpu_cpu_ic_data|altsyncram:the_altsyncram|altsyncram_ekj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 9;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 511;
defparam ram_block1a7.port_a_logical_ram_depth = 512;
defparam ram_block1a7.port_a_logical_ram_width = 32;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 9;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "none";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 511;
defparam ram_block1a7.port_b_logical_ram_depth = 512;
defparam ram_block1a7.port_b_logical_ram_width = 32;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";

cyclonev_ram_block ram_block1a20(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a20_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a20.clk0_core_clock_enable = "ena0";
defparam ram_block1a20.clk1_core_clock_enable = "ena1";
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_ic_data_module:first_nios2_system_cpu_cpu_ic_data|altsyncram:the_altsyncram|altsyncram_ekj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a20.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a20.operation_mode = "dual_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 9;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 511;
defparam ram_block1a20.port_a_logical_ram_depth = 512;
defparam ram_block1a20.port_a_logical_ram_width = 32;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a20.port_b_address_clear = "none";
defparam ram_block1a20.port_b_address_clock = "clock1";
defparam ram_block1a20.port_b_address_width = 9;
defparam ram_block1a20.port_b_data_out_clear = "none";
defparam ram_block1a20.port_b_data_out_clock = "none";
defparam ram_block1a20.port_b_data_width = 1;
defparam ram_block1a20.port_b_first_address = 0;
defparam ram_block1a20.port_b_first_bit_number = 20;
defparam ram_block1a20.port_b_last_address = 511;
defparam ram_block1a20.port_b_logical_ram_depth = 512;
defparam ram_block1a20.port_b_logical_ram_width = 32;
defparam ram_block1a20.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a20.port_b_read_enable_clock = "clock1";
defparam ram_block1a20.ram_block_type = "auto";

cyclonev_ram_block ram_block1a19(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a19_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a19.clk0_core_clock_enable = "ena0";
defparam ram_block1a19.clk1_core_clock_enable = "ena1";
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_ic_data_module:first_nios2_system_cpu_cpu_ic_data|altsyncram:the_altsyncram|altsyncram_ekj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a19.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a19.operation_mode = "dual_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 9;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 511;
defparam ram_block1a19.port_a_logical_ram_depth = 512;
defparam ram_block1a19.port_a_logical_ram_width = 32;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a19.port_b_address_clear = "none";
defparam ram_block1a19.port_b_address_clock = "clock1";
defparam ram_block1a19.port_b_address_width = 9;
defparam ram_block1a19.port_b_data_out_clear = "none";
defparam ram_block1a19.port_b_data_out_clock = "none";
defparam ram_block1a19.port_b_data_width = 1;
defparam ram_block1a19.port_b_first_address = 0;
defparam ram_block1a19.port_b_first_bit_number = 19;
defparam ram_block1a19.port_b_last_address = 511;
defparam ram_block1a19.port_b_logical_ram_depth = 512;
defparam ram_block1a19.port_b_logical_ram_width = 32;
defparam ram_block1a19.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a19.port_b_read_enable_clock = "clock1";
defparam ram_block1a19.ram_block_type = "auto";

endmodule

module first_nios2_system_first_nios2_system_cpu_cpu_ic_tag_module (
	q_b_5,
	q_b_0,
	q_b_1,
	q_b_2,
	q_b_3,
	q_b_4,
	q_b_11,
	q_b_13,
	q_b_10,
	q_b_12,
	ic_tag_wraddress_0,
	ic_tag_wraddress_1,
	ic_tag_wraddress_2,
	ic_tag_wraddress_3,
	ic_tag_wraddress_4,
	ic_tag_wraddress_5,
	ic_fill_valid_bits_5,
	ic_fill_valid_bits_7,
	ic_fill_valid_bits_4,
	q_b_7,
	q_b_9,
	q_b_6,
	q_b_8,
	ic_fill_valid_bits_6,
	ic_fill_valid_bits_1,
	ic_fill_valid_bits_3,
	ic_fill_valid_bits_0,
	ic_fill_valid_bits_2,
	ic_fill_tag_5,
	ic_fill_tag_4,
	ic_fill_tag_3,
	ic_fill_tag_2,
	ic_fill_tag_1,
	ic_fill_tag_0,
	F_stall,
	F_ic_tag_rd_addr_nxt_0,
	F_ic_tag_rd_addr_nxt_1,
	F_ic_tag_rd_addr_nxt_2,
	F_ic_tag_rd_addr_nxt_3,
	F_ic_tag_rd_addr_nxt_4,
	F_ic_tag_rd_addr_nxt_5,
	ic_tag_wren,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_5;
output 	q_b_0;
output 	q_b_1;
output 	q_b_2;
output 	q_b_3;
output 	q_b_4;
output 	q_b_11;
output 	q_b_13;
output 	q_b_10;
output 	q_b_12;
input 	ic_tag_wraddress_0;
input 	ic_tag_wraddress_1;
input 	ic_tag_wraddress_2;
input 	ic_tag_wraddress_3;
input 	ic_tag_wraddress_4;
input 	ic_tag_wraddress_5;
input 	ic_fill_valid_bits_5;
input 	ic_fill_valid_bits_7;
input 	ic_fill_valid_bits_4;
output 	q_b_7;
output 	q_b_9;
output 	q_b_6;
output 	q_b_8;
input 	ic_fill_valid_bits_6;
input 	ic_fill_valid_bits_1;
input 	ic_fill_valid_bits_3;
input 	ic_fill_valid_bits_0;
input 	ic_fill_valid_bits_2;
input 	ic_fill_tag_5;
input 	ic_fill_tag_4;
input 	ic_fill_tag_3;
input 	ic_fill_tag_2;
input 	ic_fill_tag_1;
input 	ic_fill_tag_0;
input 	F_stall;
input 	F_ic_tag_rd_addr_nxt_0;
input 	F_ic_tag_rd_addr_nxt_1;
input 	F_ic_tag_rd_addr_nxt_2;
input 	F_ic_tag_rd_addr_nxt_3;
input 	F_ic_tag_rd_addr_nxt_4;
input 	F_ic_tag_rd_addr_nxt_5;
input 	ic_tag_wren;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



first_nios2_system_altsyncram_3 the_altsyncram(
	.q_b({q_b_unconnected_wire_31,q_b_unconnected_wire_30,q_b_unconnected_wire_29,q_b_unconnected_wire_28,q_b_unconnected_wire_27,q_b_unconnected_wire_26,q_b_unconnected_wire_25,q_b_unconnected_wire_24,q_b_unconnected_wire_23,q_b_unconnected_wire_22,q_b_unconnected_wire_21,
q_b_unconnected_wire_20,q_b_unconnected_wire_19,q_b_unconnected_wire_18,q_b_unconnected_wire_17,q_b_unconnected_wire_16,q_b_unconnected_wire_15,q_b_unconnected_wire_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.address_a({gnd,gnd,gnd,gnd,gnd,gnd,gnd,ic_tag_wraddress_5,ic_tag_wraddress_4,ic_tag_wraddress_3,ic_tag_wraddress_2,ic_tag_wraddress_1,ic_tag_wraddress_0}),
	.data_a({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,ic_fill_valid_bits_7,ic_fill_valid_bits_6,ic_fill_valid_bits_5,ic_fill_valid_bits_4,ic_fill_valid_bits_3,ic_fill_valid_bits_2,ic_fill_valid_bits_1,ic_fill_valid_bits_0,ic_fill_tag_5,ic_fill_tag_4,ic_fill_tag_3,
ic_fill_tag_2,ic_fill_tag_1,ic_fill_tag_0}),
	.rden_b(F_stall),
	.address_b({gnd,gnd,gnd,F_ic_tag_rd_addr_nxt_5,F_ic_tag_rd_addr_nxt_4,F_ic_tag_rd_addr_nxt_3,F_ic_tag_rd_addr_nxt_2,F_ic_tag_rd_addr_nxt_1,F_ic_tag_rd_addr_nxt_0}),
	.wren_a(ic_tag_wren),
	.clock0(clk_clk));

endmodule

module first_nios2_system_altsyncram_3 (
	q_b,
	address_a,
	data_a,
	rden_b,
	address_b,
	wren_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_b;
input 	[12:0] address_a;
input 	[31:0] data_a;
input 	rden_b;
input 	[8:0] address_b;
input 	wren_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



first_nios2_system_altsyncram_ldj1 auto_generated(
	.q_b({q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.address_a({address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.data_a({data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.rden_b(rden_b),
	.address_b({address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.wren_a(wren_a),
	.clock0(clock0));

endmodule

module first_nios2_system_altsyncram_ldj1 (
	q_b,
	address_a,
	data_a,
	rden_b,
	address_b,
	wren_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[13:0] q_b;
input 	[5:0] address_a;
input 	[13:0] data_a;
input 	rden_b;
input 	[5:0] address_b;
input 	wren_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

cyclonev_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(!rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_ic_tag_module:first_nios2_system_cpu_cpu_ic_tag|altsyncram:the_altsyncram|altsyncram_ldj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "old";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 6;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 63;
defparam ram_block1a5.port_a_logical_ram_depth = 64;
defparam ram_block1a5.port_a_logical_ram_width = 14;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock0";
defparam ram_block1a5.port_b_address_width = 6;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "none";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 63;
defparam ram_block1a5.port_b_logical_ram_depth = 64;
defparam ram_block1a5.port_b_logical_ram_width = 14;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock0";
defparam ram_block1a5.ram_block_type = "auto";

cyclonev_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(!rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_ic_tag_module:first_nios2_system_cpu_cpu_ic_tag|altsyncram:the_altsyncram|altsyncram_ldj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "old";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 6;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 63;
defparam ram_block1a0.port_a_logical_ram_depth = 64;
defparam ram_block1a0.port_a_logical_ram_width = 14;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock0";
defparam ram_block1a0.port_b_address_width = 6;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "none";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 63;
defparam ram_block1a0.port_b_logical_ram_depth = 64;
defparam ram_block1a0.port_b_logical_ram_width = 14;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock0";
defparam ram_block1a0.ram_block_type = "auto";

cyclonev_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(!rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_ic_tag_module:first_nios2_system_cpu_cpu_ic_tag|altsyncram:the_altsyncram|altsyncram_ldj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "old";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 6;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 63;
defparam ram_block1a1.port_a_logical_ram_depth = 64;
defparam ram_block1a1.port_a_logical_ram_width = 14;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock0";
defparam ram_block1a1.port_b_address_width = 6;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "none";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 63;
defparam ram_block1a1.port_b_logical_ram_depth = 64;
defparam ram_block1a1.port_b_logical_ram_width = 14;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock0";
defparam ram_block1a1.ram_block_type = "auto";

cyclonev_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(!rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_ic_tag_module:first_nios2_system_cpu_cpu_ic_tag|altsyncram:the_altsyncram|altsyncram_ldj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "old";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 6;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 63;
defparam ram_block1a2.port_a_logical_ram_depth = 64;
defparam ram_block1a2.port_a_logical_ram_width = 14;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock0";
defparam ram_block1a2.port_b_address_width = 6;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "none";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 63;
defparam ram_block1a2.port_b_logical_ram_depth = 64;
defparam ram_block1a2.port_b_logical_ram_width = 14;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock0";
defparam ram_block1a2.ram_block_type = "auto";

cyclonev_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(!rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_ic_tag_module:first_nios2_system_cpu_cpu_ic_tag|altsyncram:the_altsyncram|altsyncram_ldj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "old";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 6;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 63;
defparam ram_block1a3.port_a_logical_ram_depth = 64;
defparam ram_block1a3.port_a_logical_ram_width = 14;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock0";
defparam ram_block1a3.port_b_address_width = 6;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "none";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 63;
defparam ram_block1a3.port_b_logical_ram_depth = 64;
defparam ram_block1a3.port_b_logical_ram_width = 14;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock0";
defparam ram_block1a3.ram_block_type = "auto";

cyclonev_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(!rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_ic_tag_module:first_nios2_system_cpu_cpu_ic_tag|altsyncram:the_altsyncram|altsyncram_ldj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "old";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 6;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 63;
defparam ram_block1a4.port_a_logical_ram_depth = 64;
defparam ram_block1a4.port_a_logical_ram_width = 14;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock0";
defparam ram_block1a4.port_b_address_width = 6;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "none";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 63;
defparam ram_block1a4.port_b_logical_ram_depth = 64;
defparam ram_block1a4.port_b_logical_ram_width = 14;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock0";
defparam ram_block1a4.ram_block_type = "auto";

cyclonev_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(!rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_ic_tag_module:first_nios2_system_cpu_cpu_ic_tag|altsyncram:the_altsyncram|altsyncram_ldj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "old";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 6;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 63;
defparam ram_block1a11.port_a_logical_ram_depth = 64;
defparam ram_block1a11.port_a_logical_ram_width = 14;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock0";
defparam ram_block1a11.port_b_address_width = 6;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "none";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 63;
defparam ram_block1a11.port_b_logical_ram_depth = 64;
defparam ram_block1a11.port_b_logical_ram_width = 14;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock0";
defparam ram_block1a11.ram_block_type = "auto";

cyclonev_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(!rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_ic_tag_module:first_nios2_system_cpu_cpu_ic_tag|altsyncram:the_altsyncram|altsyncram_ldj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "old";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 6;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 63;
defparam ram_block1a13.port_a_logical_ram_depth = 64;
defparam ram_block1a13.port_a_logical_ram_width = 14;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock0";
defparam ram_block1a13.port_b_address_width = 6;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "none";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 63;
defparam ram_block1a13.port_b_logical_ram_depth = 64;
defparam ram_block1a13.port_b_logical_ram_width = 14;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock0";
defparam ram_block1a13.ram_block_type = "auto";

cyclonev_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(!rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_ic_tag_module:first_nios2_system_cpu_cpu_ic_tag|altsyncram:the_altsyncram|altsyncram_ldj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "old";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 6;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 63;
defparam ram_block1a10.port_a_logical_ram_depth = 64;
defparam ram_block1a10.port_a_logical_ram_width = 14;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock0";
defparam ram_block1a10.port_b_address_width = 6;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "none";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 63;
defparam ram_block1a10.port_b_logical_ram_depth = 64;
defparam ram_block1a10.port_b_logical_ram_width = 14;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock0";
defparam ram_block1a10.ram_block_type = "auto";

cyclonev_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(!rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_ic_tag_module:first_nios2_system_cpu_cpu_ic_tag|altsyncram:the_altsyncram|altsyncram_ldj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "old";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 6;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 63;
defparam ram_block1a12.port_a_logical_ram_depth = 64;
defparam ram_block1a12.port_a_logical_ram_width = 14;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock0";
defparam ram_block1a12.port_b_address_width = 6;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "none";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 63;
defparam ram_block1a12.port_b_logical_ram_depth = 64;
defparam ram_block1a12.port_b_logical_ram_width = 14;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock0";
defparam ram_block1a12.ram_block_type = "auto";

cyclonev_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(!rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_ic_tag_module:first_nios2_system_cpu_cpu_ic_tag|altsyncram:the_altsyncram|altsyncram_ldj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "old";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 6;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 63;
defparam ram_block1a7.port_a_logical_ram_depth = 64;
defparam ram_block1a7.port_a_logical_ram_width = 14;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock0";
defparam ram_block1a7.port_b_address_width = 6;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "none";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 63;
defparam ram_block1a7.port_b_logical_ram_depth = 64;
defparam ram_block1a7.port_b_logical_ram_width = 14;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock0";
defparam ram_block1a7.ram_block_type = "auto";

cyclonev_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(!rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_ic_tag_module:first_nios2_system_cpu_cpu_ic_tag|altsyncram:the_altsyncram|altsyncram_ldj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "old";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 6;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 63;
defparam ram_block1a9.port_a_logical_ram_depth = 64;
defparam ram_block1a9.port_a_logical_ram_width = 14;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock0";
defparam ram_block1a9.port_b_address_width = 6;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "none";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 63;
defparam ram_block1a9.port_b_logical_ram_depth = 64;
defparam ram_block1a9.port_b_logical_ram_width = 14;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock0";
defparam ram_block1a9.ram_block_type = "auto";

cyclonev_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(!rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_ic_tag_module:first_nios2_system_cpu_cpu_ic_tag|altsyncram:the_altsyncram|altsyncram_ldj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "old";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 6;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 63;
defparam ram_block1a6.port_a_logical_ram_depth = 64;
defparam ram_block1a6.port_a_logical_ram_width = 14;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock0";
defparam ram_block1a6.port_b_address_width = 6;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "none";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 63;
defparam ram_block1a6.port_b_logical_ram_depth = 64;
defparam ram_block1a6.port_b_logical_ram_width = 14;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock0";
defparam ram_block1a6.ram_block_type = "auto";

cyclonev_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(!rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_ic_tag_module:first_nios2_system_cpu_cpu_ic_tag|altsyncram:the_altsyncram|altsyncram_ldj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "old";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 6;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 63;
defparam ram_block1a8.port_a_logical_ram_depth = 64;
defparam ram_block1a8.port_a_logical_ram_width = 14;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock0";
defparam ram_block1a8.port_b_address_width = 6;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "none";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 63;
defparam ram_block1a8.port_b_logical_ram_depth = 64;
defparam ram_block1a8.port_b_logical_ram_width = 14;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock0";
defparam ram_block1a8.ram_block_type = "auto";

endmodule

module first_nios2_system_first_nios2_system_cpu_cpu_mult_cell (
	E_src1_3,
	E_src2_22,
	E_src1_22,
	E_src2_23,
	E_src1_23,
	E_src2_24,
	E_src1_24,
	E_src1_0,
	E_src2_25,
	E_src1_25,
	E_src1_2,
	E_src1_31,
	E_src2_7,
	E_src1_7,
	E_src2_21,
	E_src1_21,
	E_src2_11,
	E_src1_11,
	E_src2_28,
	E_src1_28,
	E_src2_10,
	E_src1_10,
	E_src2_27,
	E_src1_27,
	E_src2_8,
	E_src1_8,
	E_src2_9,
	E_src1_9,
	E_src1_4,
	E_src2_5,
	E_src1_5,
	E_src2_6,
	E_src1_6,
	E_src2_26,
	E_src1_26,
	E_src2_20,
	E_src1_20,
	E_src2_19,
	E_src1_19,
	E_src2_17,
	E_src1_17,
	E_src2_30,
	E_src1_30,
	E_src1_1,
	E_src2_18,
	E_src1_18,
	E_src2_16,
	E_src1_16,
	E_src2_15,
	E_src1_15,
	E_src2_12,
	E_src1_12,
	E_src2_13,
	E_src1_13,
	E_src2_14,
	E_src1_14,
	E_src2_29,
	E_src1_29,
	r_sync_rst,
	A_mem_stall,
	E_src2_3,
	E_src2_0,
	E_src2_2,
	E_src2_31,
	E_src2_4,
	E_src2_1,
	data_out_wire_0,
	data_out_wire_1,
	data_out_wire_2,
	data_out_wire_3,
	data_out_wire_4,
	data_out_wire_5,
	data_out_wire_6,
	data_out_wire_7,
	data_out_wire_11,
	data_out_wire_10,
	data_out_wire_8,
	data_out_wire_9,
	data_out_wire_15,
	data_out_wire_12,
	data_out_wire_13,
	data_out_wire_14,
	data_out_wire_61,
	data_out_wire_71,
	data_out_wire_81,
	data_out_wire_91,
	data_out_wire_151,
	data_out_wire_51,
	data_out_wire_121,
	data_out_wire_111,
	data_out_wire_101,
	data_out_wire_41,
	data_out_wire_31,
	data_out_wire_16,
	data_out_wire_141,
	data_out_wire_21,
	data_out_wire_01,
	data_out_wire_131,
	data_out_wire_62,
	data_out_wire_22,
	data_out_wire_72,
	data_out_wire_23,
	data_out_wire_82,
	data_out_wire_24,
	data_out_wire_92,
	data_out_wire_25,
	data_out_wire_152,
	data_out_wire_311,
	data_out_wire_52,
	data_out_wire_211,
	data_out_wire_122,
	data_out_wire_28,
	data_out_wire_112,
	data_out_wire_27,
	data_out_wire_102,
	data_out_wire_26,
	data_out_wire_42,
	data_out_wire_20,
	data_out_wire_32,
	data_out_wire_19,
	data_out_wire_17,
	data_out_wire_171,
	data_out_wire_142,
	data_out_wire_30,
	data_out_wire_29,
	data_out_wire_18,
	data_out_wire_02,
	data_out_wire_161,
	data_out_wire_132,
	data_out_wire_291,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	E_src1_3;
input 	E_src2_22;
input 	E_src1_22;
input 	E_src2_23;
input 	E_src1_23;
input 	E_src2_24;
input 	E_src1_24;
input 	E_src1_0;
input 	E_src2_25;
input 	E_src1_25;
input 	E_src1_2;
input 	E_src1_31;
input 	E_src2_7;
input 	E_src1_7;
input 	E_src2_21;
input 	E_src1_21;
input 	E_src2_11;
input 	E_src1_11;
input 	E_src2_28;
input 	E_src1_28;
input 	E_src2_10;
input 	E_src1_10;
input 	E_src2_27;
input 	E_src1_27;
input 	E_src2_8;
input 	E_src1_8;
input 	E_src2_9;
input 	E_src1_9;
input 	E_src1_4;
input 	E_src2_5;
input 	E_src1_5;
input 	E_src2_6;
input 	E_src1_6;
input 	E_src2_26;
input 	E_src1_26;
input 	E_src2_20;
input 	E_src1_20;
input 	E_src2_19;
input 	E_src1_19;
input 	E_src2_17;
input 	E_src1_17;
input 	E_src2_30;
input 	E_src1_30;
input 	E_src1_1;
input 	E_src2_18;
input 	E_src1_18;
input 	E_src2_16;
input 	E_src1_16;
input 	E_src2_15;
input 	E_src1_15;
input 	E_src2_12;
input 	E_src1_12;
input 	E_src2_13;
input 	E_src1_13;
input 	E_src2_14;
input 	E_src1_14;
input 	E_src2_29;
input 	E_src1_29;
input 	r_sync_rst;
input 	A_mem_stall;
input 	E_src2_3;
input 	E_src2_0;
input 	E_src2_2;
input 	E_src2_31;
input 	E_src2_4;
input 	E_src2_1;
output 	data_out_wire_0;
output 	data_out_wire_1;
output 	data_out_wire_2;
output 	data_out_wire_3;
output 	data_out_wire_4;
output 	data_out_wire_5;
output 	data_out_wire_6;
output 	data_out_wire_7;
output 	data_out_wire_11;
output 	data_out_wire_10;
output 	data_out_wire_8;
output 	data_out_wire_9;
output 	data_out_wire_15;
output 	data_out_wire_12;
output 	data_out_wire_13;
output 	data_out_wire_14;
output 	data_out_wire_61;
output 	data_out_wire_71;
output 	data_out_wire_81;
output 	data_out_wire_91;
output 	data_out_wire_151;
output 	data_out_wire_51;
output 	data_out_wire_121;
output 	data_out_wire_111;
output 	data_out_wire_101;
output 	data_out_wire_41;
output 	data_out_wire_31;
output 	data_out_wire_16;
output 	data_out_wire_141;
output 	data_out_wire_21;
output 	data_out_wire_01;
output 	data_out_wire_131;
output 	data_out_wire_62;
output 	data_out_wire_22;
output 	data_out_wire_72;
output 	data_out_wire_23;
output 	data_out_wire_82;
output 	data_out_wire_24;
output 	data_out_wire_92;
output 	data_out_wire_25;
output 	data_out_wire_152;
output 	data_out_wire_311;
output 	data_out_wire_52;
output 	data_out_wire_211;
output 	data_out_wire_122;
output 	data_out_wire_28;
output 	data_out_wire_112;
output 	data_out_wire_27;
output 	data_out_wire_102;
output 	data_out_wire_26;
output 	data_out_wire_42;
output 	data_out_wire_20;
output 	data_out_wire_32;
output 	data_out_wire_19;
output 	data_out_wire_17;
output 	data_out_wire_171;
output 	data_out_wire_142;
output 	data_out_wire_30;
output 	data_out_wire_29;
output 	data_out_wire_18;
output 	data_out_wire_02;
output 	data_out_wire_161;
output 	data_out_wire_132;
output 	data_out_wire_291;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



first_nios2_system_altera_mult_add the_altmult_add_p1(
	.E_src1_3(E_src1_3),
	.E_src1_0(E_src1_0),
	.E_src1_2(E_src1_2),
	.E_src2_7(E_src2_7),
	.E_src1_7(E_src1_7),
	.E_src2_11(E_src2_11),
	.E_src1_11(E_src1_11),
	.E_src2_10(E_src2_10),
	.E_src1_10(E_src1_10),
	.E_src2_8(E_src2_8),
	.E_src1_8(E_src1_8),
	.E_src2_9(E_src2_9),
	.E_src1_9(E_src1_9),
	.E_src1_4(E_src1_4),
	.E_src2_5(E_src2_5),
	.E_src1_5(E_src1_5),
	.E_src2_6(E_src2_6),
	.E_src1_6(E_src1_6),
	.E_src1_1(E_src1_1),
	.E_src2_15(E_src2_15),
	.E_src1_15(E_src1_15),
	.E_src2_12(E_src2_12),
	.E_src1_12(E_src1_12),
	.E_src2_13(E_src2_13),
	.E_src1_13(E_src1_13),
	.E_src2_14(E_src2_14),
	.E_src1_14(E_src1_14),
	.r_sync_rst(r_sync_rst),
	.A_mem_stall(A_mem_stall),
	.E_src2_3(E_src2_3),
	.E_src2_0(E_src2_0),
	.E_src2_2(E_src2_2),
	.E_src2_4(E_src2_4),
	.E_src2_1(E_src2_1),
	.data_out_wire_0(data_out_wire_0),
	.data_out_wire_1(data_out_wire_1),
	.data_out_wire_2(data_out_wire_2),
	.data_out_wire_3(data_out_wire_3),
	.data_out_wire_4(data_out_wire_4),
	.data_out_wire_5(data_out_wire_5),
	.data_out_wire_6(data_out_wire_6),
	.data_out_wire_7(data_out_wire_7),
	.data_out_wire_11(data_out_wire_11),
	.data_out_wire_10(data_out_wire_10),
	.data_out_wire_8(data_out_wire_8),
	.data_out_wire_9(data_out_wire_9),
	.data_out_wire_15(data_out_wire_15),
	.data_out_wire_12(data_out_wire_12),
	.data_out_wire_13(data_out_wire_13),
	.data_out_wire_14(data_out_wire_14),
	.data_out_wire_22(data_out_wire_22),
	.data_out_wire_23(data_out_wire_23),
	.data_out_wire_24(data_out_wire_24),
	.data_out_wire_25(data_out_wire_25),
	.data_out_wire_31(data_out_wire_311),
	.data_out_wire_21(data_out_wire_211),
	.data_out_wire_28(data_out_wire_28),
	.data_out_wire_27(data_out_wire_27),
	.data_out_wire_26(data_out_wire_26),
	.data_out_wire_20(data_out_wire_20),
	.data_out_wire_19(data_out_wire_19),
	.data_out_wire_17(data_out_wire_171),
	.data_out_wire_30(data_out_wire_30),
	.data_out_wire_18(data_out_wire_18),
	.data_out_wire_16(data_out_wire_161),
	.data_out_wire_29(data_out_wire_291),
	.clk_clk(clk_clk));

first_nios2_system_altera_mult_add_2 the_altmult_add_p3(
	.E_src1_22(E_src1_22),
	.E_src1_23(E_src1_23),
	.E_src1_24(E_src1_24),
	.E_src1_25(E_src1_25),
	.E_src1_31(E_src1_31),
	.E_src2_7(E_src2_7),
	.E_src1_21(E_src1_21),
	.E_src2_11(E_src2_11),
	.E_src1_28(E_src1_28),
	.E_src2_10(E_src2_10),
	.E_src1_27(E_src1_27),
	.E_src2_8(E_src2_8),
	.E_src2_9(E_src2_9),
	.E_src2_5(E_src2_5),
	.E_src2_6(E_src2_6),
	.E_src1_26(E_src1_26),
	.E_src1_20(E_src1_20),
	.E_src1_19(E_src1_19),
	.E_src1_17(E_src1_17),
	.E_src1_30(E_src1_30),
	.E_src1_18(E_src1_18),
	.E_src1_16(E_src1_16),
	.E_src2_15(E_src2_15),
	.E_src2_12(E_src2_12),
	.E_src2_13(E_src2_13),
	.E_src2_14(E_src2_14),
	.E_src1_29(E_src1_29),
	.r_sync_rst(r_sync_rst),
	.A_mem_stall(A_mem_stall),
	.E_src2_3(E_src2_3),
	.E_src2_0(E_src2_0),
	.E_src2_2(E_src2_2),
	.E_src2_4(E_src2_4),
	.E_src2_1(E_src2_1),
	.data_out_wire_6(data_out_wire_61),
	.data_out_wire_7(data_out_wire_71),
	.data_out_wire_8(data_out_wire_81),
	.data_out_wire_9(data_out_wire_91),
	.data_out_wire_15(data_out_wire_151),
	.data_out_wire_5(data_out_wire_51),
	.data_out_wire_12(data_out_wire_121),
	.data_out_wire_11(data_out_wire_111),
	.data_out_wire_10(data_out_wire_101),
	.data_out_wire_4(data_out_wire_41),
	.data_out_wire_3(data_out_wire_31),
	.data_out_wire_1(data_out_wire_16),
	.data_out_wire_14(data_out_wire_141),
	.data_out_wire_2(data_out_wire_21),
	.data_out_wire_0(data_out_wire_01),
	.data_out_wire_13(data_out_wire_131),
	.clk_clk(clk_clk));

first_nios2_system_altera_mult_add_1 the_altmult_add_p2(
	.E_src1_3(E_src1_3),
	.E_src2_22(E_src2_22),
	.E_src2_23(E_src2_23),
	.E_src2_24(E_src2_24),
	.E_src1_0(E_src1_0),
	.E_src2_25(E_src2_25),
	.E_src1_2(E_src1_2),
	.E_src1_7(E_src1_7),
	.E_src2_21(E_src2_21),
	.E_src1_11(E_src1_11),
	.E_src2_28(E_src2_28),
	.E_src1_10(E_src1_10),
	.E_src2_27(E_src2_27),
	.E_src1_8(E_src1_8),
	.E_src1_9(E_src1_9),
	.E_src1_4(E_src1_4),
	.E_src1_5(E_src1_5),
	.E_src1_6(E_src1_6),
	.E_src2_26(E_src2_26),
	.E_src2_20(E_src2_20),
	.E_src2_19(E_src2_19),
	.E_src2_17(E_src2_17),
	.E_src2_30(E_src2_30),
	.E_src1_1(E_src1_1),
	.E_src2_18(E_src2_18),
	.E_src2_16(E_src2_16),
	.E_src1_15(E_src1_15),
	.E_src1_12(E_src1_12),
	.E_src1_13(E_src1_13),
	.E_src1_14(E_src1_14),
	.E_src2_29(E_src2_29),
	.r_sync_rst(r_sync_rst),
	.A_mem_stall(A_mem_stall),
	.E_src2_31(E_src2_31),
	.data_out_wire_6(data_out_wire_62),
	.data_out_wire_7(data_out_wire_72),
	.data_out_wire_8(data_out_wire_82),
	.data_out_wire_9(data_out_wire_92),
	.data_out_wire_15(data_out_wire_152),
	.data_out_wire_5(data_out_wire_52),
	.data_out_wire_12(data_out_wire_122),
	.data_out_wire_11(data_out_wire_112),
	.data_out_wire_10(data_out_wire_102),
	.data_out_wire_4(data_out_wire_42),
	.data_out_wire_3(data_out_wire_32),
	.data_out_wire_1(data_out_wire_17),
	.data_out_wire_14(data_out_wire_142),
	.data_out_wire_2(data_out_wire_29),
	.data_out_wire_0(data_out_wire_02),
	.data_out_wire_13(data_out_wire_132),
	.clk_clk(clk_clk));

endmodule

module first_nios2_system_altera_mult_add (
	E_src1_3,
	E_src1_0,
	E_src1_2,
	E_src2_7,
	E_src1_7,
	E_src2_11,
	E_src1_11,
	E_src2_10,
	E_src1_10,
	E_src2_8,
	E_src1_8,
	E_src2_9,
	E_src1_9,
	E_src1_4,
	E_src2_5,
	E_src1_5,
	E_src2_6,
	E_src1_6,
	E_src1_1,
	E_src2_15,
	E_src1_15,
	E_src2_12,
	E_src1_12,
	E_src2_13,
	E_src1_13,
	E_src2_14,
	E_src1_14,
	r_sync_rst,
	A_mem_stall,
	E_src2_3,
	E_src2_0,
	E_src2_2,
	E_src2_4,
	E_src2_1,
	data_out_wire_0,
	data_out_wire_1,
	data_out_wire_2,
	data_out_wire_3,
	data_out_wire_4,
	data_out_wire_5,
	data_out_wire_6,
	data_out_wire_7,
	data_out_wire_11,
	data_out_wire_10,
	data_out_wire_8,
	data_out_wire_9,
	data_out_wire_15,
	data_out_wire_12,
	data_out_wire_13,
	data_out_wire_14,
	data_out_wire_22,
	data_out_wire_23,
	data_out_wire_24,
	data_out_wire_25,
	data_out_wire_31,
	data_out_wire_21,
	data_out_wire_28,
	data_out_wire_27,
	data_out_wire_26,
	data_out_wire_20,
	data_out_wire_19,
	data_out_wire_17,
	data_out_wire_30,
	data_out_wire_18,
	data_out_wire_16,
	data_out_wire_29,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	E_src1_3;
input 	E_src1_0;
input 	E_src1_2;
input 	E_src2_7;
input 	E_src1_7;
input 	E_src2_11;
input 	E_src1_11;
input 	E_src2_10;
input 	E_src1_10;
input 	E_src2_8;
input 	E_src1_8;
input 	E_src2_9;
input 	E_src1_9;
input 	E_src1_4;
input 	E_src2_5;
input 	E_src1_5;
input 	E_src2_6;
input 	E_src1_6;
input 	E_src1_1;
input 	E_src2_15;
input 	E_src1_15;
input 	E_src2_12;
input 	E_src1_12;
input 	E_src2_13;
input 	E_src1_13;
input 	E_src2_14;
input 	E_src1_14;
input 	r_sync_rst;
input 	A_mem_stall;
input 	E_src2_3;
input 	E_src2_0;
input 	E_src2_2;
input 	E_src2_4;
input 	E_src2_1;
output 	data_out_wire_0;
output 	data_out_wire_1;
output 	data_out_wire_2;
output 	data_out_wire_3;
output 	data_out_wire_4;
output 	data_out_wire_5;
output 	data_out_wire_6;
output 	data_out_wire_7;
output 	data_out_wire_11;
output 	data_out_wire_10;
output 	data_out_wire_8;
output 	data_out_wire_9;
output 	data_out_wire_15;
output 	data_out_wire_12;
output 	data_out_wire_13;
output 	data_out_wire_14;
output 	data_out_wire_22;
output 	data_out_wire_23;
output 	data_out_wire_24;
output 	data_out_wire_25;
output 	data_out_wire_31;
output 	data_out_wire_21;
output 	data_out_wire_28;
output 	data_out_wire_27;
output 	data_out_wire_26;
output 	data_out_wire_20;
output 	data_out_wire_19;
output 	data_out_wire_17;
output 	data_out_wire_30;
output 	data_out_wire_18;
output 	data_out_wire_16;
output 	data_out_wire_29;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



first_nios2_system_altera_mult_add_37p2 auto_generated(
	.E_src1_3(E_src1_3),
	.E_src1_0(E_src1_0),
	.E_src1_2(E_src1_2),
	.E_src2_7(E_src2_7),
	.E_src1_7(E_src1_7),
	.E_src2_11(E_src2_11),
	.E_src1_11(E_src1_11),
	.E_src2_10(E_src2_10),
	.E_src1_10(E_src1_10),
	.E_src2_8(E_src2_8),
	.E_src1_8(E_src1_8),
	.E_src2_9(E_src2_9),
	.E_src1_9(E_src1_9),
	.E_src1_4(E_src1_4),
	.E_src2_5(E_src2_5),
	.E_src1_5(E_src1_5),
	.E_src2_6(E_src2_6),
	.E_src1_6(E_src1_6),
	.E_src1_1(E_src1_1),
	.E_src2_15(E_src2_15),
	.E_src1_15(E_src1_15),
	.E_src2_12(E_src2_12),
	.E_src1_12(E_src1_12),
	.E_src2_13(E_src2_13),
	.E_src1_13(E_src1_13),
	.E_src2_14(E_src2_14),
	.E_src1_14(E_src1_14),
	.r_sync_rst(r_sync_rst),
	.A_mem_stall(A_mem_stall),
	.E_src2_3(E_src2_3),
	.E_src2_0(E_src2_0),
	.E_src2_2(E_src2_2),
	.E_src2_4(E_src2_4),
	.E_src2_1(E_src2_1),
	.data_out_wire_0(data_out_wire_0),
	.data_out_wire_1(data_out_wire_1),
	.data_out_wire_2(data_out_wire_2),
	.data_out_wire_3(data_out_wire_3),
	.data_out_wire_4(data_out_wire_4),
	.data_out_wire_5(data_out_wire_5),
	.data_out_wire_6(data_out_wire_6),
	.data_out_wire_7(data_out_wire_7),
	.data_out_wire_11(data_out_wire_11),
	.data_out_wire_10(data_out_wire_10),
	.data_out_wire_8(data_out_wire_8),
	.data_out_wire_9(data_out_wire_9),
	.data_out_wire_15(data_out_wire_15),
	.data_out_wire_12(data_out_wire_12),
	.data_out_wire_13(data_out_wire_13),
	.data_out_wire_14(data_out_wire_14),
	.data_out_wire_22(data_out_wire_22),
	.data_out_wire_23(data_out_wire_23),
	.data_out_wire_24(data_out_wire_24),
	.data_out_wire_25(data_out_wire_25),
	.data_out_wire_31(data_out_wire_31),
	.data_out_wire_21(data_out_wire_21),
	.data_out_wire_28(data_out_wire_28),
	.data_out_wire_27(data_out_wire_27),
	.data_out_wire_26(data_out_wire_26),
	.data_out_wire_20(data_out_wire_20),
	.data_out_wire_19(data_out_wire_19),
	.data_out_wire_17(data_out_wire_17),
	.data_out_wire_30(data_out_wire_30),
	.data_out_wire_18(data_out_wire_18),
	.data_out_wire_16(data_out_wire_16),
	.data_out_wire_29(data_out_wire_29),
	.clk_clk(clk_clk));

endmodule

module first_nios2_system_altera_mult_add_37p2 (
	E_src1_3,
	E_src1_0,
	E_src1_2,
	E_src2_7,
	E_src1_7,
	E_src2_11,
	E_src1_11,
	E_src2_10,
	E_src1_10,
	E_src2_8,
	E_src1_8,
	E_src2_9,
	E_src1_9,
	E_src1_4,
	E_src2_5,
	E_src1_5,
	E_src2_6,
	E_src1_6,
	E_src1_1,
	E_src2_15,
	E_src1_15,
	E_src2_12,
	E_src1_12,
	E_src2_13,
	E_src1_13,
	E_src2_14,
	E_src1_14,
	r_sync_rst,
	A_mem_stall,
	E_src2_3,
	E_src2_0,
	E_src2_2,
	E_src2_4,
	E_src2_1,
	data_out_wire_0,
	data_out_wire_1,
	data_out_wire_2,
	data_out_wire_3,
	data_out_wire_4,
	data_out_wire_5,
	data_out_wire_6,
	data_out_wire_7,
	data_out_wire_11,
	data_out_wire_10,
	data_out_wire_8,
	data_out_wire_9,
	data_out_wire_15,
	data_out_wire_12,
	data_out_wire_13,
	data_out_wire_14,
	data_out_wire_22,
	data_out_wire_23,
	data_out_wire_24,
	data_out_wire_25,
	data_out_wire_31,
	data_out_wire_21,
	data_out_wire_28,
	data_out_wire_27,
	data_out_wire_26,
	data_out_wire_20,
	data_out_wire_19,
	data_out_wire_17,
	data_out_wire_30,
	data_out_wire_18,
	data_out_wire_16,
	data_out_wire_29,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	E_src1_3;
input 	E_src1_0;
input 	E_src1_2;
input 	E_src2_7;
input 	E_src1_7;
input 	E_src2_11;
input 	E_src1_11;
input 	E_src2_10;
input 	E_src1_10;
input 	E_src2_8;
input 	E_src1_8;
input 	E_src2_9;
input 	E_src1_9;
input 	E_src1_4;
input 	E_src2_5;
input 	E_src1_5;
input 	E_src2_6;
input 	E_src1_6;
input 	E_src1_1;
input 	E_src2_15;
input 	E_src1_15;
input 	E_src2_12;
input 	E_src1_12;
input 	E_src2_13;
input 	E_src1_13;
input 	E_src2_14;
input 	E_src1_14;
input 	r_sync_rst;
input 	A_mem_stall;
input 	E_src2_3;
input 	E_src2_0;
input 	E_src2_2;
input 	E_src2_4;
input 	E_src2_1;
output 	data_out_wire_0;
output 	data_out_wire_1;
output 	data_out_wire_2;
output 	data_out_wire_3;
output 	data_out_wire_4;
output 	data_out_wire_5;
output 	data_out_wire_6;
output 	data_out_wire_7;
output 	data_out_wire_11;
output 	data_out_wire_10;
output 	data_out_wire_8;
output 	data_out_wire_9;
output 	data_out_wire_15;
output 	data_out_wire_12;
output 	data_out_wire_13;
output 	data_out_wire_14;
output 	data_out_wire_22;
output 	data_out_wire_23;
output 	data_out_wire_24;
output 	data_out_wire_25;
output 	data_out_wire_31;
output 	data_out_wire_21;
output 	data_out_wire_28;
output 	data_out_wire_27;
output 	data_out_wire_26;
output 	data_out_wire_20;
output 	data_out_wire_19;
output 	data_out_wire_17;
output 	data_out_wire_30;
output 	data_out_wire_18;
output 	data_out_wire_16;
output 	data_out_wire_29;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



first_nios2_system_altera_mult_add_rtl_1 altera_mult_add_rtl1(
	.E_src1_3(E_src1_3),
	.E_src1_0(E_src1_0),
	.E_src1_2(E_src1_2),
	.E_src2_7(E_src2_7),
	.E_src1_7(E_src1_7),
	.E_src2_11(E_src2_11),
	.E_src1_11(E_src1_11),
	.E_src2_10(E_src2_10),
	.E_src1_10(E_src1_10),
	.E_src2_8(E_src2_8),
	.E_src1_8(E_src1_8),
	.E_src2_9(E_src2_9),
	.E_src1_9(E_src1_9),
	.E_src1_4(E_src1_4),
	.E_src2_5(E_src2_5),
	.E_src1_5(E_src1_5),
	.E_src2_6(E_src2_6),
	.E_src1_6(E_src1_6),
	.E_src1_1(E_src1_1),
	.E_src2_15(E_src2_15),
	.E_src1_15(E_src1_15),
	.E_src2_12(E_src2_12),
	.E_src1_12(E_src1_12),
	.E_src2_13(E_src2_13),
	.E_src1_13(E_src1_13),
	.E_src2_14(E_src2_14),
	.E_src1_14(E_src1_14),
	.r_sync_rst(r_sync_rst),
	.A_mem_stall(A_mem_stall),
	.E_src2_3(E_src2_3),
	.E_src2_0(E_src2_0),
	.E_src2_2(E_src2_2),
	.E_src2_4(E_src2_4),
	.E_src2_1(E_src2_1),
	.data_out_wire_0(data_out_wire_0),
	.data_out_wire_1(data_out_wire_1),
	.data_out_wire_2(data_out_wire_2),
	.data_out_wire_3(data_out_wire_3),
	.data_out_wire_4(data_out_wire_4),
	.data_out_wire_5(data_out_wire_5),
	.data_out_wire_6(data_out_wire_6),
	.data_out_wire_7(data_out_wire_7),
	.data_out_wire_11(data_out_wire_11),
	.data_out_wire_10(data_out_wire_10),
	.data_out_wire_8(data_out_wire_8),
	.data_out_wire_9(data_out_wire_9),
	.data_out_wire_15(data_out_wire_15),
	.data_out_wire_12(data_out_wire_12),
	.data_out_wire_13(data_out_wire_13),
	.data_out_wire_14(data_out_wire_14),
	.data_out_wire_22(data_out_wire_22),
	.data_out_wire_23(data_out_wire_23),
	.data_out_wire_24(data_out_wire_24),
	.data_out_wire_25(data_out_wire_25),
	.data_out_wire_31(data_out_wire_31),
	.data_out_wire_21(data_out_wire_21),
	.data_out_wire_28(data_out_wire_28),
	.data_out_wire_27(data_out_wire_27),
	.data_out_wire_26(data_out_wire_26),
	.data_out_wire_20(data_out_wire_20),
	.data_out_wire_19(data_out_wire_19),
	.data_out_wire_17(data_out_wire_17),
	.data_out_wire_30(data_out_wire_30),
	.data_out_wire_18(data_out_wire_18),
	.data_out_wire_16(data_out_wire_16),
	.data_out_wire_29(data_out_wire_29),
	.clk_clk(clk_clk));

endmodule

module first_nios2_system_altera_mult_add_rtl_1 (
	E_src1_3,
	E_src1_0,
	E_src1_2,
	E_src2_7,
	E_src1_7,
	E_src2_11,
	E_src1_11,
	E_src2_10,
	E_src1_10,
	E_src2_8,
	E_src1_8,
	E_src2_9,
	E_src1_9,
	E_src1_4,
	E_src2_5,
	E_src1_5,
	E_src2_6,
	E_src1_6,
	E_src1_1,
	E_src2_15,
	E_src1_15,
	E_src2_12,
	E_src1_12,
	E_src2_13,
	E_src1_13,
	E_src2_14,
	E_src1_14,
	r_sync_rst,
	A_mem_stall,
	E_src2_3,
	E_src2_0,
	E_src2_2,
	E_src2_4,
	E_src2_1,
	data_out_wire_0,
	data_out_wire_1,
	data_out_wire_2,
	data_out_wire_3,
	data_out_wire_4,
	data_out_wire_5,
	data_out_wire_6,
	data_out_wire_7,
	data_out_wire_11,
	data_out_wire_10,
	data_out_wire_8,
	data_out_wire_9,
	data_out_wire_15,
	data_out_wire_12,
	data_out_wire_13,
	data_out_wire_14,
	data_out_wire_22,
	data_out_wire_23,
	data_out_wire_24,
	data_out_wire_25,
	data_out_wire_31,
	data_out_wire_21,
	data_out_wire_28,
	data_out_wire_27,
	data_out_wire_26,
	data_out_wire_20,
	data_out_wire_19,
	data_out_wire_17,
	data_out_wire_30,
	data_out_wire_18,
	data_out_wire_16,
	data_out_wire_29,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	E_src1_3;
input 	E_src1_0;
input 	E_src1_2;
input 	E_src2_7;
input 	E_src1_7;
input 	E_src2_11;
input 	E_src1_11;
input 	E_src2_10;
input 	E_src1_10;
input 	E_src2_8;
input 	E_src1_8;
input 	E_src2_9;
input 	E_src1_9;
input 	E_src1_4;
input 	E_src2_5;
input 	E_src1_5;
input 	E_src2_6;
input 	E_src1_6;
input 	E_src1_1;
input 	E_src2_15;
input 	E_src1_15;
input 	E_src2_12;
input 	E_src1_12;
input 	E_src2_13;
input 	E_src1_13;
input 	E_src2_14;
input 	E_src1_14;
input 	r_sync_rst;
input 	A_mem_stall;
input 	E_src2_3;
input 	E_src2_0;
input 	E_src2_2;
input 	E_src2_4;
input 	E_src2_1;
output 	data_out_wire_0;
output 	data_out_wire_1;
output 	data_out_wire_2;
output 	data_out_wire_3;
output 	data_out_wire_4;
output 	data_out_wire_5;
output 	data_out_wire_6;
output 	data_out_wire_7;
output 	data_out_wire_11;
output 	data_out_wire_10;
output 	data_out_wire_8;
output 	data_out_wire_9;
output 	data_out_wire_15;
output 	data_out_wire_12;
output 	data_out_wire_13;
output 	data_out_wire_14;
output 	data_out_wire_22;
output 	data_out_wire_23;
output 	data_out_wire_24;
output 	data_out_wire_25;
output 	data_out_wire_31;
output 	data_out_wire_21;
output 	data_out_wire_28;
output 	data_out_wire_27;
output 	data_out_wire_26;
output 	data_out_wire_20;
output 	data_out_wire_19;
output 	data_out_wire_17;
output 	data_out_wire_30;
output 	data_out_wire_18;
output 	data_out_wire_16;
output 	data_out_wire_29;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



first_nios2_system_ama_multiplier_function multiplier_block(
	.E_src1_3(E_src1_3),
	.E_src1_0(E_src1_0),
	.E_src1_2(E_src1_2),
	.E_src2_7(E_src2_7),
	.E_src1_7(E_src1_7),
	.E_src2_11(E_src2_11),
	.E_src1_11(E_src1_11),
	.E_src2_10(E_src2_10),
	.E_src1_10(E_src1_10),
	.E_src2_8(E_src2_8),
	.E_src1_8(E_src1_8),
	.E_src2_9(E_src2_9),
	.E_src1_9(E_src1_9),
	.E_src1_4(E_src1_4),
	.E_src2_5(E_src2_5),
	.E_src1_5(E_src1_5),
	.E_src2_6(E_src2_6),
	.E_src1_6(E_src1_6),
	.E_src1_1(E_src1_1),
	.E_src2_15(E_src2_15),
	.E_src1_15(E_src1_15),
	.E_src2_12(E_src2_12),
	.E_src1_12(E_src1_12),
	.E_src2_13(E_src2_13),
	.E_src1_13(E_src1_13),
	.E_src2_14(E_src2_14),
	.E_src1_14(E_src1_14),
	.r_sync_rst(r_sync_rst),
	.A_mem_stall(A_mem_stall),
	.E_src2_3(E_src2_3),
	.E_src2_0(E_src2_0),
	.E_src2_2(E_src2_2),
	.E_src2_4(E_src2_4),
	.E_src2_1(E_src2_1),
	.data_out_wire_0(data_out_wire_0),
	.data_out_wire_1(data_out_wire_1),
	.data_out_wire_2(data_out_wire_2),
	.data_out_wire_3(data_out_wire_3),
	.data_out_wire_4(data_out_wire_4),
	.data_out_wire_5(data_out_wire_5),
	.data_out_wire_6(data_out_wire_6),
	.data_out_wire_7(data_out_wire_7),
	.data_out_wire_11(data_out_wire_11),
	.data_out_wire_10(data_out_wire_10),
	.data_out_wire_8(data_out_wire_8),
	.data_out_wire_9(data_out_wire_9),
	.data_out_wire_15(data_out_wire_15),
	.data_out_wire_12(data_out_wire_12),
	.data_out_wire_13(data_out_wire_13),
	.data_out_wire_14(data_out_wire_14),
	.data_out_wire_22(data_out_wire_22),
	.data_out_wire_23(data_out_wire_23),
	.data_out_wire_24(data_out_wire_24),
	.data_out_wire_25(data_out_wire_25),
	.data_out_wire_31(data_out_wire_31),
	.data_out_wire_21(data_out_wire_21),
	.data_out_wire_28(data_out_wire_28),
	.data_out_wire_27(data_out_wire_27),
	.data_out_wire_26(data_out_wire_26),
	.data_out_wire_20(data_out_wire_20),
	.data_out_wire_19(data_out_wire_19),
	.data_out_wire_17(data_out_wire_17),
	.data_out_wire_30(data_out_wire_30),
	.data_out_wire_18(data_out_wire_18),
	.data_out_wire_16(data_out_wire_16),
	.data_out_wire_29(data_out_wire_29),
	.clk_clk(clk_clk));

endmodule

module first_nios2_system_ama_multiplier_function (
	E_src1_3,
	E_src1_0,
	E_src1_2,
	E_src2_7,
	E_src1_7,
	E_src2_11,
	E_src1_11,
	E_src2_10,
	E_src1_10,
	E_src2_8,
	E_src1_8,
	E_src2_9,
	E_src1_9,
	E_src1_4,
	E_src2_5,
	E_src1_5,
	E_src2_6,
	E_src1_6,
	E_src1_1,
	E_src2_15,
	E_src1_15,
	E_src2_12,
	E_src1_12,
	E_src2_13,
	E_src1_13,
	E_src2_14,
	E_src1_14,
	r_sync_rst,
	A_mem_stall,
	E_src2_3,
	E_src2_0,
	E_src2_2,
	E_src2_4,
	E_src2_1,
	data_out_wire_0,
	data_out_wire_1,
	data_out_wire_2,
	data_out_wire_3,
	data_out_wire_4,
	data_out_wire_5,
	data_out_wire_6,
	data_out_wire_7,
	data_out_wire_11,
	data_out_wire_10,
	data_out_wire_8,
	data_out_wire_9,
	data_out_wire_15,
	data_out_wire_12,
	data_out_wire_13,
	data_out_wire_14,
	data_out_wire_22,
	data_out_wire_23,
	data_out_wire_24,
	data_out_wire_25,
	data_out_wire_31,
	data_out_wire_21,
	data_out_wire_28,
	data_out_wire_27,
	data_out_wire_26,
	data_out_wire_20,
	data_out_wire_19,
	data_out_wire_17,
	data_out_wire_30,
	data_out_wire_18,
	data_out_wire_16,
	data_out_wire_29,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	E_src1_3;
input 	E_src1_0;
input 	E_src1_2;
input 	E_src2_7;
input 	E_src1_7;
input 	E_src2_11;
input 	E_src1_11;
input 	E_src2_10;
input 	E_src1_10;
input 	E_src2_8;
input 	E_src1_8;
input 	E_src2_9;
input 	E_src1_9;
input 	E_src1_4;
input 	E_src2_5;
input 	E_src1_5;
input 	E_src2_6;
input 	E_src1_6;
input 	E_src1_1;
input 	E_src2_15;
input 	E_src1_15;
input 	E_src2_12;
input 	E_src1_12;
input 	E_src2_13;
input 	E_src1_13;
input 	E_src2_14;
input 	E_src1_14;
input 	r_sync_rst;
input 	A_mem_stall;
input 	E_src2_3;
input 	E_src2_0;
input 	E_src2_2;
input 	E_src2_4;
input 	E_src2_1;
output 	data_out_wire_0;
output 	data_out_wire_1;
output 	data_out_wire_2;
output 	data_out_wire_3;
output 	data_out_wire_4;
output 	data_out_wire_5;
output 	data_out_wire_6;
output 	data_out_wire_7;
output 	data_out_wire_11;
output 	data_out_wire_10;
output 	data_out_wire_8;
output 	data_out_wire_9;
output 	data_out_wire_15;
output 	data_out_wire_12;
output 	data_out_wire_13;
output 	data_out_wire_14;
output 	data_out_wire_22;
output 	data_out_wire_23;
output 	data_out_wire_24;
output 	data_out_wire_25;
output 	data_out_wire_31;
output 	data_out_wire_21;
output 	data_out_wire_28;
output 	data_out_wire_27;
output 	data_out_wire_26;
output 	data_out_wire_20;
output 	data_out_wire_19;
output 	data_out_wire_17;
output 	data_out_wire_30;
output 	data_out_wire_18;
output 	data_out_wire_16;
output 	data_out_wire_29;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \data_out_wire_0[0] ;
wire \data_out_wire_0[1] ;
wire \data_out_wire_0[2] ;
wire \data_out_wire_0[3] ;
wire \data_out_wire_0[4] ;
wire \data_out_wire_0[5] ;
wire \data_out_wire_0[6] ;
wire \data_out_wire_0[7] ;
wire \data_out_wire_0[8] ;
wire \data_out_wire_0[9] ;
wire \data_out_wire_0[10] ;
wire \data_out_wire_0[11] ;
wire \data_out_wire_0[12] ;
wire \data_out_wire_0[13] ;
wire \data_out_wire_0[14] ;
wire \data_out_wire_0[15] ;
wire \data_out_wire_0[16] ;
wire \data_out_wire_0[17] ;
wire \data_out_wire_0[18] ;
wire \data_out_wire_0[19] ;
wire \data_out_wire_0[20] ;
wire \data_out_wire_0[21] ;
wire \data_out_wire_0[22] ;
wire \data_out_wire_0[23] ;
wire \data_out_wire_0[24] ;
wire \data_out_wire_0[25] ;
wire \data_out_wire_0[26] ;
wire \data_out_wire_0[27] ;
wire \data_out_wire_0[28] ;
wire \data_out_wire_0[29] ;
wire \data_out_wire_0[30] ;
wire \data_out_wire_0[31] ;
wire \Mult0~8 ;
wire \Mult0~9 ;
wire \Mult0~10 ;
wire \Mult0~11 ;
wire \Mult0~12 ;
wire \Mult0~13 ;
wire \Mult0~14 ;
wire \Mult0~15 ;
wire \Mult0~16 ;
wire \Mult0~17 ;
wire \Mult0~18 ;
wire \Mult0~19 ;
wire \Mult0~20 ;
wire \Mult0~21 ;
wire \Mult0~22 ;
wire \Mult0~23 ;
wire \Mult0~24 ;
wire \Mult0~25 ;
wire \Mult0~26 ;
wire \Mult0~27 ;
wire \Mult0~28 ;
wire \Mult0~29 ;
wire \Mult0~30 ;
wire \Mult0~31 ;
wire \Mult0~32 ;
wire \Mult0~33 ;
wire \Mult0~34 ;
wire \Mult0~35 ;
wire \Mult0~36 ;
wire \Mult0~37 ;
wire \Mult0~38 ;
wire \Mult0~39 ;

wire [63:0] \Mult0~mac_RESULTA_bus ;

assign \data_out_wire_0[0]  = \Mult0~mac_RESULTA_bus [0];
assign \data_out_wire_0[1]  = \Mult0~mac_RESULTA_bus [1];
assign \data_out_wire_0[2]  = \Mult0~mac_RESULTA_bus [2];
assign \data_out_wire_0[3]  = \Mult0~mac_RESULTA_bus [3];
assign \data_out_wire_0[4]  = \Mult0~mac_RESULTA_bus [4];
assign \data_out_wire_0[5]  = \Mult0~mac_RESULTA_bus [5];
assign \data_out_wire_0[6]  = \Mult0~mac_RESULTA_bus [6];
assign \data_out_wire_0[7]  = \Mult0~mac_RESULTA_bus [7];
assign \data_out_wire_0[8]  = \Mult0~mac_RESULTA_bus [8];
assign \data_out_wire_0[9]  = \Mult0~mac_RESULTA_bus [9];
assign \data_out_wire_0[10]  = \Mult0~mac_RESULTA_bus [10];
assign \data_out_wire_0[11]  = \Mult0~mac_RESULTA_bus [11];
assign \data_out_wire_0[12]  = \Mult0~mac_RESULTA_bus [12];
assign \data_out_wire_0[13]  = \Mult0~mac_RESULTA_bus [13];
assign \data_out_wire_0[14]  = \Mult0~mac_RESULTA_bus [14];
assign \data_out_wire_0[15]  = \Mult0~mac_RESULTA_bus [15];
assign \data_out_wire_0[16]  = \Mult0~mac_RESULTA_bus [16];
assign \data_out_wire_0[17]  = \Mult0~mac_RESULTA_bus [17];
assign \data_out_wire_0[18]  = \Mult0~mac_RESULTA_bus [18];
assign \data_out_wire_0[19]  = \Mult0~mac_RESULTA_bus [19];
assign \data_out_wire_0[20]  = \Mult0~mac_RESULTA_bus [20];
assign \data_out_wire_0[21]  = \Mult0~mac_RESULTA_bus [21];
assign \data_out_wire_0[22]  = \Mult0~mac_RESULTA_bus [22];
assign \data_out_wire_0[23]  = \Mult0~mac_RESULTA_bus [23];
assign \data_out_wire_0[24]  = \Mult0~mac_RESULTA_bus [24];
assign \data_out_wire_0[25]  = \Mult0~mac_RESULTA_bus [25];
assign \data_out_wire_0[26]  = \Mult0~mac_RESULTA_bus [26];
assign \data_out_wire_0[27]  = \Mult0~mac_RESULTA_bus [27];
assign \data_out_wire_0[28]  = \Mult0~mac_RESULTA_bus [28];
assign \data_out_wire_0[29]  = \Mult0~mac_RESULTA_bus [29];
assign \data_out_wire_0[30]  = \Mult0~mac_RESULTA_bus [30];
assign \data_out_wire_0[31]  = \Mult0~mac_RESULTA_bus [31];
assign \Mult0~8  = \Mult0~mac_RESULTA_bus [32];
assign \Mult0~9  = \Mult0~mac_RESULTA_bus [33];
assign \Mult0~10  = \Mult0~mac_RESULTA_bus [34];
assign \Mult0~11  = \Mult0~mac_RESULTA_bus [35];
assign \Mult0~12  = \Mult0~mac_RESULTA_bus [36];
assign \Mult0~13  = \Mult0~mac_RESULTA_bus [37];
assign \Mult0~14  = \Mult0~mac_RESULTA_bus [38];
assign \Mult0~15  = \Mult0~mac_RESULTA_bus [39];
assign \Mult0~16  = \Mult0~mac_RESULTA_bus [40];
assign \Mult0~17  = \Mult0~mac_RESULTA_bus [41];
assign \Mult0~18  = \Mult0~mac_RESULTA_bus [42];
assign \Mult0~19  = \Mult0~mac_RESULTA_bus [43];
assign \Mult0~20  = \Mult0~mac_RESULTA_bus [44];
assign \Mult0~21  = \Mult0~mac_RESULTA_bus [45];
assign \Mult0~22  = \Mult0~mac_RESULTA_bus [46];
assign \Mult0~23  = \Mult0~mac_RESULTA_bus [47];
assign \Mult0~24  = \Mult0~mac_RESULTA_bus [48];
assign \Mult0~25  = \Mult0~mac_RESULTA_bus [49];
assign \Mult0~26  = \Mult0~mac_RESULTA_bus [50];
assign \Mult0~27  = \Mult0~mac_RESULTA_bus [51];
assign \Mult0~28  = \Mult0~mac_RESULTA_bus [52];
assign \Mult0~29  = \Mult0~mac_RESULTA_bus [53];
assign \Mult0~30  = \Mult0~mac_RESULTA_bus [54];
assign \Mult0~31  = \Mult0~mac_RESULTA_bus [55];
assign \Mult0~32  = \Mult0~mac_RESULTA_bus [56];
assign \Mult0~33  = \Mult0~mac_RESULTA_bus [57];
assign \Mult0~34  = \Mult0~mac_RESULTA_bus [58];
assign \Mult0~35  = \Mult0~mac_RESULTA_bus [59];
assign \Mult0~36  = \Mult0~mac_RESULTA_bus [60];
assign \Mult0~37  = \Mult0~mac_RESULTA_bus [61];
assign \Mult0~38  = \Mult0~mac_RESULTA_bus [62];
assign \Mult0~39  = \Mult0~mac_RESULTA_bus [63];

first_nios2_system_ama_register_function_12 multiplier_register_block_0(
	.data_in({gnd,gnd,\data_out_wire_0[31] ,\data_out_wire_0[30] ,\data_out_wire_0[29] ,\data_out_wire_0[28] ,\data_out_wire_0[27] ,\data_out_wire_0[26] ,\data_out_wire_0[25] ,\data_out_wire_0[24] ,\data_out_wire_0[23] ,\data_out_wire_0[22] ,\data_out_wire_0[21] ,
\data_out_wire_0[20] ,\data_out_wire_0[19] ,\data_out_wire_0[18] ,\data_out_wire_0[17] ,\data_out_wire_0[16] ,\data_out_wire_0[15] ,\data_out_wire_0[14] ,\data_out_wire_0[13] ,\data_out_wire_0[12] ,\data_out_wire_0[11] ,\data_out_wire_0[10] ,\data_out_wire_0[9] ,
\data_out_wire_0[8] ,\data_out_wire_0[7] ,\data_out_wire_0[6] ,\data_out_wire_0[5] ,\data_out_wire_0[4] ,\data_out_wire_0[3] ,\data_out_wire_0[2] ,\data_out_wire_0[1] ,\data_out_wire_0[0] }),
	.aclr({gnd,gnd,gnd,r_sync_rst}),
	.ena({gnd,gnd,gnd,A_mem_stall}),
	.data_out_wire_0(data_out_wire_0),
	.data_out_wire_1(data_out_wire_1),
	.data_out_wire_2(data_out_wire_2),
	.data_out_wire_3(data_out_wire_3),
	.data_out_wire_4(data_out_wire_4),
	.data_out_wire_5(data_out_wire_5),
	.data_out_wire_6(data_out_wire_6),
	.data_out_wire_7(data_out_wire_7),
	.data_out_wire_11(data_out_wire_11),
	.data_out_wire_10(data_out_wire_10),
	.data_out_wire_8(data_out_wire_8),
	.data_out_wire_9(data_out_wire_9),
	.data_out_wire_15(data_out_wire_15),
	.data_out_wire_12(data_out_wire_12),
	.data_out_wire_13(data_out_wire_13),
	.data_out_wire_14(data_out_wire_14),
	.data_out_wire_22(data_out_wire_22),
	.data_out_wire_23(data_out_wire_23),
	.data_out_wire_24(data_out_wire_24),
	.data_out_wire_25(data_out_wire_25),
	.data_out_wire_31(data_out_wire_31),
	.data_out_wire_21(data_out_wire_21),
	.data_out_wire_28(data_out_wire_28),
	.data_out_wire_27(data_out_wire_27),
	.data_out_wire_26(data_out_wire_26),
	.data_out_wire_20(data_out_wire_20),
	.data_out_wire_19(data_out_wire_19),
	.data_out_wire_17(data_out_wire_17),
	.data_out_wire_30(data_out_wire_30),
	.data_out_wire_18(data_out_wire_18),
	.data_out_wire_16(data_out_wire_16),
	.data_out_wire_29(data_out_wire_29),
	.clock({gnd,gnd,gnd,clk_clk}));

cyclonev_mac \Mult0~mac (
	.sub(gnd),
	.negate(gnd),
	.accumulate(gnd),
	.loadconst(gnd),
	.ax({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,E_src2_15,E_src2_14,E_src2_13,E_src2_12,E_src2_11,E_src2_10,E_src2_9,E_src2_8,E_src2_7,E_src2_6,E_src2_5,E_src2_4,E_src2_3,E_src2_2,E_src2_1,E_src2_0}),
	.ay({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,E_src1_15,E_src1_14,E_src1_13,E_src1_12,E_src1_11,E_src1_10,E_src1_9,E_src1_8,E_src1_7,E_src1_6,E_src1_5,E_src1_4,E_src1_3,E_src1_2,E_src1_1,E_src1_0}),
	.az(26'b00000000000000000000000000),
	.bx(18'b000000000000000000),
	.by(19'b0000000000000000000),
	.bz(18'b000000000000000000),
	.coefsela(3'b000),
	.coefselb(3'b000),
	.clk(3'b000),
	.aclr(2'b00),
	.ena(3'b111),
	.scanin(27'b000000000000000000000000000),
	.chainin(1'b0),
	.dftout(),
	.resulta(\Mult0~mac_RESULTA_bus ),
	.resultb(),
	.scanout(),
	.chainout());
defparam \Mult0~mac .accumulate_clock = "none";
defparam \Mult0~mac .ax_clock = "none";
defparam \Mult0~mac .ax_width = 16;
defparam \Mult0~mac .ay_scan_in_clock = "none";
defparam \Mult0~mac .ay_scan_in_width = 16;
defparam \Mult0~mac .ay_use_scan_in = "false";
defparam \Mult0~mac .az_clock = "none";
defparam \Mult0~mac .bx_clock = "none";
defparam \Mult0~mac .by_clock = "none";
defparam \Mult0~mac .by_use_scan_in = "false";
defparam \Mult0~mac .bz_clock = "none";
defparam \Mult0~mac .coef_a_0 = 0;
defparam \Mult0~mac .coef_a_1 = 0;
defparam \Mult0~mac .coef_a_2 = 0;
defparam \Mult0~mac .coef_a_3 = 0;
defparam \Mult0~mac .coef_a_4 = 0;
defparam \Mult0~mac .coef_a_5 = 0;
defparam \Mult0~mac .coef_a_6 = 0;
defparam \Mult0~mac .coef_a_7 = 0;
defparam \Mult0~mac .coef_b_0 = 0;
defparam \Mult0~mac .coef_b_1 = 0;
defparam \Mult0~mac .coef_b_2 = 0;
defparam \Mult0~mac .coef_b_3 = 0;
defparam \Mult0~mac .coef_b_4 = 0;
defparam \Mult0~mac .coef_b_5 = 0;
defparam \Mult0~mac .coef_b_6 = 0;
defparam \Mult0~mac .coef_b_7 = 0;
defparam \Mult0~mac .coef_sel_a_clock = "none";
defparam \Mult0~mac .coef_sel_b_clock = "none";
defparam \Mult0~mac .delay_scan_out_ay = "false";
defparam \Mult0~mac .delay_scan_out_by = "false";
defparam \Mult0~mac .enable_double_accum = "false";
defparam \Mult0~mac .load_const_clock = "none";
defparam \Mult0~mac .load_const_value = 0;
defparam \Mult0~mac .mode_sub_location = 0;
defparam \Mult0~mac .negate_clock = "none";
defparam \Mult0~mac .operand_source_max = "input";
defparam \Mult0~mac .operand_source_may = "input";
defparam \Mult0~mac .operand_source_mbx = "input";
defparam \Mult0~mac .operand_source_mby = "input";
defparam \Mult0~mac .operation_mode = "m18x18_full";
defparam \Mult0~mac .output_clock = "none";
defparam \Mult0~mac .preadder_subtract_a = "false";
defparam \Mult0~mac .preadder_subtract_b = "false";
defparam \Mult0~mac .result_a_width = 64;
defparam \Mult0~mac .signed_max = "false";
defparam \Mult0~mac .signed_may = "false";
defparam \Mult0~mac .signed_mbx = "false";
defparam \Mult0~mac .signed_mby = "false";
defparam \Mult0~mac .sub_clock = "none";
defparam \Mult0~mac .use_chainadder = "false";

endmodule

module first_nios2_system_ama_register_function_12 (
	data_in,
	aclr,
	ena,
	data_out_wire_0,
	data_out_wire_1,
	data_out_wire_2,
	data_out_wire_3,
	data_out_wire_4,
	data_out_wire_5,
	data_out_wire_6,
	data_out_wire_7,
	data_out_wire_11,
	data_out_wire_10,
	data_out_wire_8,
	data_out_wire_9,
	data_out_wire_15,
	data_out_wire_12,
	data_out_wire_13,
	data_out_wire_14,
	data_out_wire_22,
	data_out_wire_23,
	data_out_wire_24,
	data_out_wire_25,
	data_out_wire_31,
	data_out_wire_21,
	data_out_wire_28,
	data_out_wire_27,
	data_out_wire_26,
	data_out_wire_20,
	data_out_wire_19,
	data_out_wire_17,
	data_out_wire_30,
	data_out_wire_18,
	data_out_wire_16,
	data_out_wire_29,
	clock)/* synthesis synthesis_greybox=1 */;
input 	[33:0] data_in;
input 	[3:0] aclr;
input 	[3:0] ena;
output 	data_out_wire_0;
output 	data_out_wire_1;
output 	data_out_wire_2;
output 	data_out_wire_3;
output 	data_out_wire_4;
output 	data_out_wire_5;
output 	data_out_wire_6;
output 	data_out_wire_7;
output 	data_out_wire_11;
output 	data_out_wire_10;
output 	data_out_wire_8;
output 	data_out_wire_9;
output 	data_out_wire_15;
output 	data_out_wire_12;
output 	data_out_wire_13;
output 	data_out_wire_14;
output 	data_out_wire_22;
output 	data_out_wire_23;
output 	data_out_wire_24;
output 	data_out_wire_25;
output 	data_out_wire_31;
output 	data_out_wire_21;
output 	data_out_wire_28;
output 	data_out_wire_27;
output 	data_out_wire_26;
output 	data_out_wire_20;
output 	data_out_wire_19;
output 	data_out_wire_17;
output 	data_out_wire_30;
output 	data_out_wire_18;
output 	data_out_wire_16;
output 	data_out_wire_29;
input 	[3:0] clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \data_out_wire[0] (
	.clk(clock[0]),
	.d(data_in[0]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!ena[0]),
	.q(data_out_wire_0),
	.prn(vcc));
defparam \data_out_wire[0] .is_wysiwyg = "true";
defparam \data_out_wire[0] .power_up = "low";

dffeas \data_out_wire[1] (
	.clk(clock[0]),
	.d(data_in[1]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!ena[0]),
	.q(data_out_wire_1),
	.prn(vcc));
defparam \data_out_wire[1] .is_wysiwyg = "true";
defparam \data_out_wire[1] .power_up = "low";

dffeas \data_out_wire[2] (
	.clk(clock[0]),
	.d(data_in[2]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!ena[0]),
	.q(data_out_wire_2),
	.prn(vcc));
defparam \data_out_wire[2] .is_wysiwyg = "true";
defparam \data_out_wire[2] .power_up = "low";

dffeas \data_out_wire[3] (
	.clk(clock[0]),
	.d(data_in[3]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!ena[0]),
	.q(data_out_wire_3),
	.prn(vcc));
defparam \data_out_wire[3] .is_wysiwyg = "true";
defparam \data_out_wire[3] .power_up = "low";

dffeas \data_out_wire[4] (
	.clk(clock[0]),
	.d(data_in[4]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!ena[0]),
	.q(data_out_wire_4),
	.prn(vcc));
defparam \data_out_wire[4] .is_wysiwyg = "true";
defparam \data_out_wire[4] .power_up = "low";

dffeas \data_out_wire[5] (
	.clk(clock[0]),
	.d(data_in[5]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!ena[0]),
	.q(data_out_wire_5),
	.prn(vcc));
defparam \data_out_wire[5] .is_wysiwyg = "true";
defparam \data_out_wire[5] .power_up = "low";

dffeas \data_out_wire[6] (
	.clk(clock[0]),
	.d(data_in[6]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!ena[0]),
	.q(data_out_wire_6),
	.prn(vcc));
defparam \data_out_wire[6] .is_wysiwyg = "true";
defparam \data_out_wire[6] .power_up = "low";

dffeas \data_out_wire[7] (
	.clk(clock[0]),
	.d(data_in[7]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!ena[0]),
	.q(data_out_wire_7),
	.prn(vcc));
defparam \data_out_wire[7] .is_wysiwyg = "true";
defparam \data_out_wire[7] .power_up = "low";

dffeas \data_out_wire[11] (
	.clk(clock[0]),
	.d(data_in[11]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!ena[0]),
	.q(data_out_wire_11),
	.prn(vcc));
defparam \data_out_wire[11] .is_wysiwyg = "true";
defparam \data_out_wire[11] .power_up = "low";

dffeas \data_out_wire[10] (
	.clk(clock[0]),
	.d(data_in[10]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!ena[0]),
	.q(data_out_wire_10),
	.prn(vcc));
defparam \data_out_wire[10] .is_wysiwyg = "true";
defparam \data_out_wire[10] .power_up = "low";

dffeas \data_out_wire[8] (
	.clk(clock[0]),
	.d(data_in[8]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!ena[0]),
	.q(data_out_wire_8),
	.prn(vcc));
defparam \data_out_wire[8] .is_wysiwyg = "true";
defparam \data_out_wire[8] .power_up = "low";

dffeas \data_out_wire[9] (
	.clk(clock[0]),
	.d(data_in[9]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!ena[0]),
	.q(data_out_wire_9),
	.prn(vcc));
defparam \data_out_wire[9] .is_wysiwyg = "true";
defparam \data_out_wire[9] .power_up = "low";

dffeas \data_out_wire[15] (
	.clk(clock[0]),
	.d(data_in[15]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!ena[0]),
	.q(data_out_wire_15),
	.prn(vcc));
defparam \data_out_wire[15] .is_wysiwyg = "true";
defparam \data_out_wire[15] .power_up = "low";

dffeas \data_out_wire[12] (
	.clk(clock[0]),
	.d(data_in[12]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!ena[0]),
	.q(data_out_wire_12),
	.prn(vcc));
defparam \data_out_wire[12] .is_wysiwyg = "true";
defparam \data_out_wire[12] .power_up = "low";

dffeas \data_out_wire[13] (
	.clk(clock[0]),
	.d(data_in[13]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!ena[0]),
	.q(data_out_wire_13),
	.prn(vcc));
defparam \data_out_wire[13] .is_wysiwyg = "true";
defparam \data_out_wire[13] .power_up = "low";

dffeas \data_out_wire[14] (
	.clk(clock[0]),
	.d(data_in[14]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!ena[0]),
	.q(data_out_wire_14),
	.prn(vcc));
defparam \data_out_wire[14] .is_wysiwyg = "true";
defparam \data_out_wire[14] .power_up = "low";

dffeas \data_out_wire[22] (
	.clk(clock[0]),
	.d(data_in[22]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!ena[0]),
	.q(data_out_wire_22),
	.prn(vcc));
defparam \data_out_wire[22] .is_wysiwyg = "true";
defparam \data_out_wire[22] .power_up = "low";

dffeas \data_out_wire[23] (
	.clk(clock[0]),
	.d(data_in[23]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!ena[0]),
	.q(data_out_wire_23),
	.prn(vcc));
defparam \data_out_wire[23] .is_wysiwyg = "true";
defparam \data_out_wire[23] .power_up = "low";

dffeas \data_out_wire[24] (
	.clk(clock[0]),
	.d(data_in[24]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!ena[0]),
	.q(data_out_wire_24),
	.prn(vcc));
defparam \data_out_wire[24] .is_wysiwyg = "true";
defparam \data_out_wire[24] .power_up = "low";

dffeas \data_out_wire[25] (
	.clk(clock[0]),
	.d(data_in[25]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!ena[0]),
	.q(data_out_wire_25),
	.prn(vcc));
defparam \data_out_wire[25] .is_wysiwyg = "true";
defparam \data_out_wire[25] .power_up = "low";

dffeas \data_out_wire[31] (
	.clk(clock[0]),
	.d(data_in[31]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!ena[0]),
	.q(data_out_wire_31),
	.prn(vcc));
defparam \data_out_wire[31] .is_wysiwyg = "true";
defparam \data_out_wire[31] .power_up = "low";

dffeas \data_out_wire[21] (
	.clk(clock[0]),
	.d(data_in[21]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!ena[0]),
	.q(data_out_wire_21),
	.prn(vcc));
defparam \data_out_wire[21] .is_wysiwyg = "true";
defparam \data_out_wire[21] .power_up = "low";

dffeas \data_out_wire[28] (
	.clk(clock[0]),
	.d(data_in[28]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!ena[0]),
	.q(data_out_wire_28),
	.prn(vcc));
defparam \data_out_wire[28] .is_wysiwyg = "true";
defparam \data_out_wire[28] .power_up = "low";

dffeas \data_out_wire[27] (
	.clk(clock[0]),
	.d(data_in[27]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!ena[0]),
	.q(data_out_wire_27),
	.prn(vcc));
defparam \data_out_wire[27] .is_wysiwyg = "true";
defparam \data_out_wire[27] .power_up = "low";

dffeas \data_out_wire[26] (
	.clk(clock[0]),
	.d(data_in[26]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!ena[0]),
	.q(data_out_wire_26),
	.prn(vcc));
defparam \data_out_wire[26] .is_wysiwyg = "true";
defparam \data_out_wire[26] .power_up = "low";

dffeas \data_out_wire[20] (
	.clk(clock[0]),
	.d(data_in[20]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!ena[0]),
	.q(data_out_wire_20),
	.prn(vcc));
defparam \data_out_wire[20] .is_wysiwyg = "true";
defparam \data_out_wire[20] .power_up = "low";

dffeas \data_out_wire[19] (
	.clk(clock[0]),
	.d(data_in[19]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!ena[0]),
	.q(data_out_wire_19),
	.prn(vcc));
defparam \data_out_wire[19] .is_wysiwyg = "true";
defparam \data_out_wire[19] .power_up = "low";

dffeas \data_out_wire[17] (
	.clk(clock[0]),
	.d(data_in[17]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!ena[0]),
	.q(data_out_wire_17),
	.prn(vcc));
defparam \data_out_wire[17] .is_wysiwyg = "true";
defparam \data_out_wire[17] .power_up = "low";

dffeas \data_out_wire[30] (
	.clk(clock[0]),
	.d(data_in[30]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!ena[0]),
	.q(data_out_wire_30),
	.prn(vcc));
defparam \data_out_wire[30] .is_wysiwyg = "true";
defparam \data_out_wire[30] .power_up = "low";

dffeas \data_out_wire[18] (
	.clk(clock[0]),
	.d(data_in[18]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!ena[0]),
	.q(data_out_wire_18),
	.prn(vcc));
defparam \data_out_wire[18] .is_wysiwyg = "true";
defparam \data_out_wire[18] .power_up = "low";

dffeas \data_out_wire[16] (
	.clk(clock[0]),
	.d(data_in[16]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!ena[0]),
	.q(data_out_wire_16),
	.prn(vcc));
defparam \data_out_wire[16] .is_wysiwyg = "true";
defparam \data_out_wire[16] .power_up = "low";

dffeas \data_out_wire[29] (
	.clk(clock[0]),
	.d(data_in[29]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!ena[0]),
	.q(data_out_wire_29),
	.prn(vcc));
defparam \data_out_wire[29] .is_wysiwyg = "true";
defparam \data_out_wire[29] .power_up = "low";

endmodule

module first_nios2_system_altera_mult_add_1 (
	E_src1_3,
	E_src2_22,
	E_src2_23,
	E_src2_24,
	E_src1_0,
	E_src2_25,
	E_src1_2,
	E_src1_7,
	E_src2_21,
	E_src1_11,
	E_src2_28,
	E_src1_10,
	E_src2_27,
	E_src1_8,
	E_src1_9,
	E_src1_4,
	E_src1_5,
	E_src1_6,
	E_src2_26,
	E_src2_20,
	E_src2_19,
	E_src2_17,
	E_src2_30,
	E_src1_1,
	E_src2_18,
	E_src2_16,
	E_src1_15,
	E_src1_12,
	E_src1_13,
	E_src1_14,
	E_src2_29,
	r_sync_rst,
	A_mem_stall,
	E_src2_31,
	data_out_wire_6,
	data_out_wire_7,
	data_out_wire_8,
	data_out_wire_9,
	data_out_wire_15,
	data_out_wire_5,
	data_out_wire_12,
	data_out_wire_11,
	data_out_wire_10,
	data_out_wire_4,
	data_out_wire_3,
	data_out_wire_1,
	data_out_wire_14,
	data_out_wire_2,
	data_out_wire_0,
	data_out_wire_13,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	E_src1_3;
input 	E_src2_22;
input 	E_src2_23;
input 	E_src2_24;
input 	E_src1_0;
input 	E_src2_25;
input 	E_src1_2;
input 	E_src1_7;
input 	E_src2_21;
input 	E_src1_11;
input 	E_src2_28;
input 	E_src1_10;
input 	E_src2_27;
input 	E_src1_8;
input 	E_src1_9;
input 	E_src1_4;
input 	E_src1_5;
input 	E_src1_6;
input 	E_src2_26;
input 	E_src2_20;
input 	E_src2_19;
input 	E_src2_17;
input 	E_src2_30;
input 	E_src1_1;
input 	E_src2_18;
input 	E_src2_16;
input 	E_src1_15;
input 	E_src1_12;
input 	E_src1_13;
input 	E_src1_14;
input 	E_src2_29;
input 	r_sync_rst;
input 	A_mem_stall;
input 	E_src2_31;
output 	data_out_wire_6;
output 	data_out_wire_7;
output 	data_out_wire_8;
output 	data_out_wire_9;
output 	data_out_wire_15;
output 	data_out_wire_5;
output 	data_out_wire_12;
output 	data_out_wire_11;
output 	data_out_wire_10;
output 	data_out_wire_4;
output 	data_out_wire_3;
output 	data_out_wire_1;
output 	data_out_wire_14;
output 	data_out_wire_2;
output 	data_out_wire_0;
output 	data_out_wire_13;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



first_nios2_system_altera_mult_add_37p2_1 auto_generated(
	.E_src1_3(E_src1_3),
	.E_src2_22(E_src2_22),
	.E_src2_23(E_src2_23),
	.E_src2_24(E_src2_24),
	.E_src1_0(E_src1_0),
	.E_src2_25(E_src2_25),
	.E_src1_2(E_src1_2),
	.E_src1_7(E_src1_7),
	.E_src2_21(E_src2_21),
	.E_src1_11(E_src1_11),
	.E_src2_28(E_src2_28),
	.E_src1_10(E_src1_10),
	.E_src2_27(E_src2_27),
	.E_src1_8(E_src1_8),
	.E_src1_9(E_src1_9),
	.E_src1_4(E_src1_4),
	.E_src1_5(E_src1_5),
	.E_src1_6(E_src1_6),
	.E_src2_26(E_src2_26),
	.E_src2_20(E_src2_20),
	.E_src2_19(E_src2_19),
	.E_src2_17(E_src2_17),
	.E_src2_30(E_src2_30),
	.E_src1_1(E_src1_1),
	.E_src2_18(E_src2_18),
	.E_src2_16(E_src2_16),
	.E_src1_15(E_src1_15),
	.E_src1_12(E_src1_12),
	.E_src1_13(E_src1_13),
	.E_src1_14(E_src1_14),
	.E_src2_29(E_src2_29),
	.r_sync_rst(r_sync_rst),
	.A_mem_stall(A_mem_stall),
	.E_src2_31(E_src2_31),
	.data_out_wire_6(data_out_wire_6),
	.data_out_wire_7(data_out_wire_7),
	.data_out_wire_8(data_out_wire_8),
	.data_out_wire_9(data_out_wire_9),
	.data_out_wire_15(data_out_wire_15),
	.data_out_wire_5(data_out_wire_5),
	.data_out_wire_12(data_out_wire_12),
	.data_out_wire_11(data_out_wire_11),
	.data_out_wire_10(data_out_wire_10),
	.data_out_wire_4(data_out_wire_4),
	.data_out_wire_3(data_out_wire_3),
	.data_out_wire_1(data_out_wire_1),
	.data_out_wire_14(data_out_wire_14),
	.data_out_wire_2(data_out_wire_2),
	.data_out_wire_0(data_out_wire_0),
	.data_out_wire_13(data_out_wire_13),
	.clk_clk(clk_clk));

endmodule

module first_nios2_system_altera_mult_add_37p2_1 (
	E_src1_3,
	E_src2_22,
	E_src2_23,
	E_src2_24,
	E_src1_0,
	E_src2_25,
	E_src1_2,
	E_src1_7,
	E_src2_21,
	E_src1_11,
	E_src2_28,
	E_src1_10,
	E_src2_27,
	E_src1_8,
	E_src1_9,
	E_src1_4,
	E_src1_5,
	E_src1_6,
	E_src2_26,
	E_src2_20,
	E_src2_19,
	E_src2_17,
	E_src2_30,
	E_src1_1,
	E_src2_18,
	E_src2_16,
	E_src1_15,
	E_src1_12,
	E_src1_13,
	E_src1_14,
	E_src2_29,
	r_sync_rst,
	A_mem_stall,
	E_src2_31,
	data_out_wire_6,
	data_out_wire_7,
	data_out_wire_8,
	data_out_wire_9,
	data_out_wire_15,
	data_out_wire_5,
	data_out_wire_12,
	data_out_wire_11,
	data_out_wire_10,
	data_out_wire_4,
	data_out_wire_3,
	data_out_wire_1,
	data_out_wire_14,
	data_out_wire_2,
	data_out_wire_0,
	data_out_wire_13,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	E_src1_3;
input 	E_src2_22;
input 	E_src2_23;
input 	E_src2_24;
input 	E_src1_0;
input 	E_src2_25;
input 	E_src1_2;
input 	E_src1_7;
input 	E_src2_21;
input 	E_src1_11;
input 	E_src2_28;
input 	E_src1_10;
input 	E_src2_27;
input 	E_src1_8;
input 	E_src1_9;
input 	E_src1_4;
input 	E_src1_5;
input 	E_src1_6;
input 	E_src2_26;
input 	E_src2_20;
input 	E_src2_19;
input 	E_src2_17;
input 	E_src2_30;
input 	E_src1_1;
input 	E_src2_18;
input 	E_src2_16;
input 	E_src1_15;
input 	E_src1_12;
input 	E_src1_13;
input 	E_src1_14;
input 	E_src2_29;
input 	r_sync_rst;
input 	A_mem_stall;
input 	E_src2_31;
output 	data_out_wire_6;
output 	data_out_wire_7;
output 	data_out_wire_8;
output 	data_out_wire_9;
output 	data_out_wire_15;
output 	data_out_wire_5;
output 	data_out_wire_12;
output 	data_out_wire_11;
output 	data_out_wire_10;
output 	data_out_wire_4;
output 	data_out_wire_3;
output 	data_out_wire_1;
output 	data_out_wire_14;
output 	data_out_wire_2;
output 	data_out_wire_0;
output 	data_out_wire_13;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



first_nios2_system_altera_mult_add_rtl_2 altera_mult_add_rtl1(
	.E_src1_3(E_src1_3),
	.E_src2_22(E_src2_22),
	.E_src2_23(E_src2_23),
	.E_src2_24(E_src2_24),
	.E_src1_0(E_src1_0),
	.E_src2_25(E_src2_25),
	.E_src1_2(E_src1_2),
	.E_src1_7(E_src1_7),
	.E_src2_21(E_src2_21),
	.E_src1_11(E_src1_11),
	.E_src2_28(E_src2_28),
	.E_src1_10(E_src1_10),
	.E_src2_27(E_src2_27),
	.E_src1_8(E_src1_8),
	.E_src1_9(E_src1_9),
	.E_src1_4(E_src1_4),
	.E_src1_5(E_src1_5),
	.E_src1_6(E_src1_6),
	.E_src2_26(E_src2_26),
	.E_src2_20(E_src2_20),
	.E_src2_19(E_src2_19),
	.E_src2_17(E_src2_17),
	.E_src2_30(E_src2_30),
	.E_src1_1(E_src1_1),
	.E_src2_18(E_src2_18),
	.E_src2_16(E_src2_16),
	.E_src1_15(E_src1_15),
	.E_src1_12(E_src1_12),
	.E_src1_13(E_src1_13),
	.E_src1_14(E_src1_14),
	.E_src2_29(E_src2_29),
	.r_sync_rst(r_sync_rst),
	.A_mem_stall(A_mem_stall),
	.E_src2_31(E_src2_31),
	.data_out_wire_6(data_out_wire_6),
	.data_out_wire_7(data_out_wire_7),
	.data_out_wire_8(data_out_wire_8),
	.data_out_wire_9(data_out_wire_9),
	.data_out_wire_15(data_out_wire_15),
	.data_out_wire_5(data_out_wire_5),
	.data_out_wire_12(data_out_wire_12),
	.data_out_wire_11(data_out_wire_11),
	.data_out_wire_10(data_out_wire_10),
	.data_out_wire_4(data_out_wire_4),
	.data_out_wire_3(data_out_wire_3),
	.data_out_wire_1(data_out_wire_1),
	.data_out_wire_14(data_out_wire_14),
	.data_out_wire_2(data_out_wire_2),
	.data_out_wire_0(data_out_wire_0),
	.data_out_wire_13(data_out_wire_13),
	.clk_clk(clk_clk));

endmodule

module first_nios2_system_altera_mult_add_rtl_2 (
	E_src1_3,
	E_src2_22,
	E_src2_23,
	E_src2_24,
	E_src1_0,
	E_src2_25,
	E_src1_2,
	E_src1_7,
	E_src2_21,
	E_src1_11,
	E_src2_28,
	E_src1_10,
	E_src2_27,
	E_src1_8,
	E_src1_9,
	E_src1_4,
	E_src1_5,
	E_src1_6,
	E_src2_26,
	E_src2_20,
	E_src2_19,
	E_src2_17,
	E_src2_30,
	E_src1_1,
	E_src2_18,
	E_src2_16,
	E_src1_15,
	E_src1_12,
	E_src1_13,
	E_src1_14,
	E_src2_29,
	r_sync_rst,
	A_mem_stall,
	E_src2_31,
	data_out_wire_6,
	data_out_wire_7,
	data_out_wire_8,
	data_out_wire_9,
	data_out_wire_15,
	data_out_wire_5,
	data_out_wire_12,
	data_out_wire_11,
	data_out_wire_10,
	data_out_wire_4,
	data_out_wire_3,
	data_out_wire_1,
	data_out_wire_14,
	data_out_wire_2,
	data_out_wire_0,
	data_out_wire_13,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	E_src1_3;
input 	E_src2_22;
input 	E_src2_23;
input 	E_src2_24;
input 	E_src1_0;
input 	E_src2_25;
input 	E_src1_2;
input 	E_src1_7;
input 	E_src2_21;
input 	E_src1_11;
input 	E_src2_28;
input 	E_src1_10;
input 	E_src2_27;
input 	E_src1_8;
input 	E_src1_9;
input 	E_src1_4;
input 	E_src1_5;
input 	E_src1_6;
input 	E_src2_26;
input 	E_src2_20;
input 	E_src2_19;
input 	E_src2_17;
input 	E_src2_30;
input 	E_src1_1;
input 	E_src2_18;
input 	E_src2_16;
input 	E_src1_15;
input 	E_src1_12;
input 	E_src1_13;
input 	E_src1_14;
input 	E_src2_29;
input 	r_sync_rst;
input 	A_mem_stall;
input 	E_src2_31;
output 	data_out_wire_6;
output 	data_out_wire_7;
output 	data_out_wire_8;
output 	data_out_wire_9;
output 	data_out_wire_15;
output 	data_out_wire_5;
output 	data_out_wire_12;
output 	data_out_wire_11;
output 	data_out_wire_10;
output 	data_out_wire_4;
output 	data_out_wire_3;
output 	data_out_wire_1;
output 	data_out_wire_14;
output 	data_out_wire_2;
output 	data_out_wire_0;
output 	data_out_wire_13;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



first_nios2_system_ama_multiplier_function_1 multiplier_block(
	.E_src1_3(E_src1_3),
	.E_src2_22(E_src2_22),
	.E_src2_23(E_src2_23),
	.E_src2_24(E_src2_24),
	.E_src1_0(E_src1_0),
	.E_src2_25(E_src2_25),
	.E_src1_2(E_src1_2),
	.E_src1_7(E_src1_7),
	.E_src2_21(E_src2_21),
	.E_src1_11(E_src1_11),
	.E_src2_28(E_src2_28),
	.E_src1_10(E_src1_10),
	.E_src2_27(E_src2_27),
	.E_src1_8(E_src1_8),
	.E_src1_9(E_src1_9),
	.E_src1_4(E_src1_4),
	.E_src1_5(E_src1_5),
	.E_src1_6(E_src1_6),
	.E_src2_26(E_src2_26),
	.E_src2_20(E_src2_20),
	.E_src2_19(E_src2_19),
	.E_src2_17(E_src2_17),
	.E_src2_30(E_src2_30),
	.E_src1_1(E_src1_1),
	.E_src2_18(E_src2_18),
	.E_src2_16(E_src2_16),
	.E_src1_15(E_src1_15),
	.E_src1_12(E_src1_12),
	.E_src1_13(E_src1_13),
	.E_src1_14(E_src1_14),
	.E_src2_29(E_src2_29),
	.r_sync_rst(r_sync_rst),
	.A_mem_stall(A_mem_stall),
	.E_src2_31(E_src2_31),
	.data_out_wire_6(data_out_wire_6),
	.data_out_wire_7(data_out_wire_7),
	.data_out_wire_8(data_out_wire_8),
	.data_out_wire_9(data_out_wire_9),
	.data_out_wire_15(data_out_wire_15),
	.data_out_wire_5(data_out_wire_5),
	.data_out_wire_12(data_out_wire_12),
	.data_out_wire_11(data_out_wire_11),
	.data_out_wire_10(data_out_wire_10),
	.data_out_wire_4(data_out_wire_4),
	.data_out_wire_3(data_out_wire_3),
	.data_out_wire_1(data_out_wire_1),
	.data_out_wire_14(data_out_wire_14),
	.data_out_wire_2(data_out_wire_2),
	.data_out_wire_0(data_out_wire_0),
	.data_out_wire_13(data_out_wire_13),
	.clk_clk(clk_clk));

endmodule

module first_nios2_system_ama_multiplier_function_1 (
	E_src1_3,
	E_src2_22,
	E_src2_23,
	E_src2_24,
	E_src1_0,
	E_src2_25,
	E_src1_2,
	E_src1_7,
	E_src2_21,
	E_src1_11,
	E_src2_28,
	E_src1_10,
	E_src2_27,
	E_src1_8,
	E_src1_9,
	E_src1_4,
	E_src1_5,
	E_src1_6,
	E_src2_26,
	E_src2_20,
	E_src2_19,
	E_src2_17,
	E_src2_30,
	E_src1_1,
	E_src2_18,
	E_src2_16,
	E_src1_15,
	E_src1_12,
	E_src1_13,
	E_src1_14,
	E_src2_29,
	r_sync_rst,
	A_mem_stall,
	E_src2_31,
	data_out_wire_6,
	data_out_wire_7,
	data_out_wire_8,
	data_out_wire_9,
	data_out_wire_15,
	data_out_wire_5,
	data_out_wire_12,
	data_out_wire_11,
	data_out_wire_10,
	data_out_wire_4,
	data_out_wire_3,
	data_out_wire_1,
	data_out_wire_14,
	data_out_wire_2,
	data_out_wire_0,
	data_out_wire_13,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	E_src1_3;
input 	E_src2_22;
input 	E_src2_23;
input 	E_src2_24;
input 	E_src1_0;
input 	E_src2_25;
input 	E_src1_2;
input 	E_src1_7;
input 	E_src2_21;
input 	E_src1_11;
input 	E_src2_28;
input 	E_src1_10;
input 	E_src2_27;
input 	E_src1_8;
input 	E_src1_9;
input 	E_src1_4;
input 	E_src1_5;
input 	E_src1_6;
input 	E_src2_26;
input 	E_src2_20;
input 	E_src2_19;
input 	E_src2_17;
input 	E_src2_30;
input 	E_src1_1;
input 	E_src2_18;
input 	E_src2_16;
input 	E_src1_15;
input 	E_src1_12;
input 	E_src1_13;
input 	E_src1_14;
input 	E_src2_29;
input 	r_sync_rst;
input 	A_mem_stall;
input 	E_src2_31;
output 	data_out_wire_6;
output 	data_out_wire_7;
output 	data_out_wire_8;
output 	data_out_wire_9;
output 	data_out_wire_15;
output 	data_out_wire_5;
output 	data_out_wire_12;
output 	data_out_wire_11;
output 	data_out_wire_10;
output 	data_out_wire_4;
output 	data_out_wire_3;
output 	data_out_wire_1;
output 	data_out_wire_14;
output 	data_out_wire_2;
output 	data_out_wire_0;
output 	data_out_wire_13;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \data_out_wire_0[0] ;
wire \data_out_wire_0[1] ;
wire \data_out_wire_0[2] ;
wire \data_out_wire_0[3] ;
wire \data_out_wire_0[4] ;
wire \data_out_wire_0[5] ;
wire \data_out_wire_0[6] ;
wire \data_out_wire_0[7] ;
wire \data_out_wire_0[8] ;
wire \data_out_wire_0[9] ;
wire \data_out_wire_0[10] ;
wire \data_out_wire_0[11] ;
wire \data_out_wire_0[12] ;
wire \data_out_wire_0[13] ;
wire \data_out_wire_0[14] ;
wire \data_out_wire_0[15] ;
wire \Mult0~8 ;
wire \Mult0~9 ;
wire \Mult0~10 ;
wire \Mult0~11 ;
wire \Mult0~12 ;
wire \Mult0~13 ;
wire \Mult0~14 ;
wire \Mult0~15 ;
wire \Mult0~16 ;
wire \Mult0~17 ;
wire \Mult0~18 ;
wire \Mult0~19 ;
wire \Mult0~20 ;
wire \Mult0~21 ;
wire \Mult0~22 ;
wire \Mult0~23 ;
wire \Mult0~24 ;
wire \Mult0~25 ;
wire \Mult0~26 ;
wire \Mult0~27 ;
wire \Mult0~28 ;
wire \Mult0~29 ;
wire \Mult0~30 ;
wire \Mult0~31 ;
wire \Mult0~32 ;
wire \Mult0~33 ;
wire \Mult0~34 ;
wire \Mult0~35 ;
wire \Mult0~36 ;
wire \Mult0~37 ;
wire \Mult0~38 ;
wire \Mult0~39 ;
wire \Mult0~40 ;
wire \Mult0~41 ;
wire \Mult0~42 ;
wire \Mult0~43 ;
wire \Mult0~44 ;
wire \Mult0~45 ;
wire \Mult0~46 ;
wire \Mult0~47 ;
wire \Mult0~48 ;
wire \Mult0~49 ;
wire \Mult0~50 ;
wire \Mult0~51 ;
wire \Mult0~52 ;
wire \Mult0~53 ;
wire \Mult0~54 ;
wire \Mult0~55 ;

wire [63:0] \Mult0~mac_RESULTA_bus ;

assign \data_out_wire_0[0]  = \Mult0~mac_RESULTA_bus [0];
assign \data_out_wire_0[1]  = \Mult0~mac_RESULTA_bus [1];
assign \data_out_wire_0[2]  = \Mult0~mac_RESULTA_bus [2];
assign \data_out_wire_0[3]  = \Mult0~mac_RESULTA_bus [3];
assign \data_out_wire_0[4]  = \Mult0~mac_RESULTA_bus [4];
assign \data_out_wire_0[5]  = \Mult0~mac_RESULTA_bus [5];
assign \data_out_wire_0[6]  = \Mult0~mac_RESULTA_bus [6];
assign \data_out_wire_0[7]  = \Mult0~mac_RESULTA_bus [7];
assign \data_out_wire_0[8]  = \Mult0~mac_RESULTA_bus [8];
assign \data_out_wire_0[9]  = \Mult0~mac_RESULTA_bus [9];
assign \data_out_wire_0[10]  = \Mult0~mac_RESULTA_bus [10];
assign \data_out_wire_0[11]  = \Mult0~mac_RESULTA_bus [11];
assign \data_out_wire_0[12]  = \Mult0~mac_RESULTA_bus [12];
assign \data_out_wire_0[13]  = \Mult0~mac_RESULTA_bus [13];
assign \data_out_wire_0[14]  = \Mult0~mac_RESULTA_bus [14];
assign \data_out_wire_0[15]  = \Mult0~mac_RESULTA_bus [15];
assign \Mult0~8  = \Mult0~mac_RESULTA_bus [16];
assign \Mult0~9  = \Mult0~mac_RESULTA_bus [17];
assign \Mult0~10  = \Mult0~mac_RESULTA_bus [18];
assign \Mult0~11  = \Mult0~mac_RESULTA_bus [19];
assign \Mult0~12  = \Mult0~mac_RESULTA_bus [20];
assign \Mult0~13  = \Mult0~mac_RESULTA_bus [21];
assign \Mult0~14  = \Mult0~mac_RESULTA_bus [22];
assign \Mult0~15  = \Mult0~mac_RESULTA_bus [23];
assign \Mult0~16  = \Mult0~mac_RESULTA_bus [24];
assign \Mult0~17  = \Mult0~mac_RESULTA_bus [25];
assign \Mult0~18  = \Mult0~mac_RESULTA_bus [26];
assign \Mult0~19  = \Mult0~mac_RESULTA_bus [27];
assign \Mult0~20  = \Mult0~mac_RESULTA_bus [28];
assign \Mult0~21  = \Mult0~mac_RESULTA_bus [29];
assign \Mult0~22  = \Mult0~mac_RESULTA_bus [30];
assign \Mult0~23  = \Mult0~mac_RESULTA_bus [31];
assign \Mult0~24  = \Mult0~mac_RESULTA_bus [32];
assign \Mult0~25  = \Mult0~mac_RESULTA_bus [33];
assign \Mult0~26  = \Mult0~mac_RESULTA_bus [34];
assign \Mult0~27  = \Mult0~mac_RESULTA_bus [35];
assign \Mult0~28  = \Mult0~mac_RESULTA_bus [36];
assign \Mult0~29  = \Mult0~mac_RESULTA_bus [37];
assign \Mult0~30  = \Mult0~mac_RESULTA_bus [38];
assign \Mult0~31  = \Mult0~mac_RESULTA_bus [39];
assign \Mult0~32  = \Mult0~mac_RESULTA_bus [40];
assign \Mult0~33  = \Mult0~mac_RESULTA_bus [41];
assign \Mult0~34  = \Mult0~mac_RESULTA_bus [42];
assign \Mult0~35  = \Mult0~mac_RESULTA_bus [43];
assign \Mult0~36  = \Mult0~mac_RESULTA_bus [44];
assign \Mult0~37  = \Mult0~mac_RESULTA_bus [45];
assign \Mult0~38  = \Mult0~mac_RESULTA_bus [46];
assign \Mult0~39  = \Mult0~mac_RESULTA_bus [47];
assign \Mult0~40  = \Mult0~mac_RESULTA_bus [48];
assign \Mult0~41  = \Mult0~mac_RESULTA_bus [49];
assign \Mult0~42  = \Mult0~mac_RESULTA_bus [50];
assign \Mult0~43  = \Mult0~mac_RESULTA_bus [51];
assign \Mult0~44  = \Mult0~mac_RESULTA_bus [52];
assign \Mult0~45  = \Mult0~mac_RESULTA_bus [53];
assign \Mult0~46  = \Mult0~mac_RESULTA_bus [54];
assign \Mult0~47  = \Mult0~mac_RESULTA_bus [55];
assign \Mult0~48  = \Mult0~mac_RESULTA_bus [56];
assign \Mult0~49  = \Mult0~mac_RESULTA_bus [57];
assign \Mult0~50  = \Mult0~mac_RESULTA_bus [58];
assign \Mult0~51  = \Mult0~mac_RESULTA_bus [59];
assign \Mult0~52  = \Mult0~mac_RESULTA_bus [60];
assign \Mult0~53  = \Mult0~mac_RESULTA_bus [61];
assign \Mult0~54  = \Mult0~mac_RESULTA_bus [62];
assign \Mult0~55  = \Mult0~mac_RESULTA_bus [63];

first_nios2_system_ama_register_function_31 multiplier_register_block_0(
	.data_in({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\data_out_wire_0[15] ,\data_out_wire_0[14] ,\data_out_wire_0[13] ,\data_out_wire_0[12] ,\data_out_wire_0[11] ,\data_out_wire_0[10] ,\data_out_wire_0[9] ,\data_out_wire_0[8] ,\data_out_wire_0[7] ,
\data_out_wire_0[6] ,\data_out_wire_0[5] ,\data_out_wire_0[4] ,\data_out_wire_0[3] ,\data_out_wire_0[2] ,\data_out_wire_0[1] ,\data_out_wire_0[0] }),
	.aclr({gnd,gnd,gnd,r_sync_rst}),
	.ena({gnd,gnd,gnd,A_mem_stall}),
	.data_out_wire_6(data_out_wire_6),
	.data_out_wire_7(data_out_wire_7),
	.data_out_wire_8(data_out_wire_8),
	.data_out_wire_9(data_out_wire_9),
	.data_out_wire_15(data_out_wire_15),
	.data_out_wire_5(data_out_wire_5),
	.data_out_wire_12(data_out_wire_12),
	.data_out_wire_11(data_out_wire_11),
	.data_out_wire_10(data_out_wire_10),
	.data_out_wire_4(data_out_wire_4),
	.data_out_wire_3(data_out_wire_3),
	.data_out_wire_1(data_out_wire_1),
	.data_out_wire_14(data_out_wire_14),
	.data_out_wire_2(data_out_wire_2),
	.data_out_wire_0(data_out_wire_0),
	.data_out_wire_13(data_out_wire_13),
	.clock({gnd,gnd,gnd,clk_clk}));

cyclonev_mac \Mult0~mac (
	.sub(gnd),
	.negate(gnd),
	.accumulate(gnd),
	.loadconst(gnd),
	.ax({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,E_src2_31,E_src2_30,E_src2_29,E_src2_28,E_src2_27,E_src2_26,E_src2_25,E_src2_24,E_src2_23,E_src2_22,E_src2_21,E_src2_20,E_src2_19,E_src2_18,E_src2_17,E_src2_16}),
	.ay({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,E_src1_15,E_src1_14,E_src1_13,E_src1_12,E_src1_11,E_src1_10,E_src1_9,E_src1_8,E_src1_7,E_src1_6,E_src1_5,E_src1_4,E_src1_3,E_src1_2,E_src1_1,E_src1_0}),
	.az(26'b00000000000000000000000000),
	.bx(18'b000000000000000000),
	.by(19'b0000000000000000000),
	.bz(18'b000000000000000000),
	.coefsela(3'b000),
	.coefselb(3'b000),
	.clk(3'b000),
	.aclr(2'b00),
	.ena(3'b111),
	.scanin(27'b000000000000000000000000000),
	.chainin(1'b0),
	.dftout(),
	.resulta(\Mult0~mac_RESULTA_bus ),
	.resultb(),
	.scanout(),
	.chainout());
defparam \Mult0~mac .accumulate_clock = "none";
defparam \Mult0~mac .ax_clock = "none";
defparam \Mult0~mac .ax_width = 16;
defparam \Mult0~mac .ay_scan_in_clock = "none";
defparam \Mult0~mac .ay_scan_in_width = 16;
defparam \Mult0~mac .ay_use_scan_in = "false";
defparam \Mult0~mac .az_clock = "none";
defparam \Mult0~mac .bx_clock = "none";
defparam \Mult0~mac .by_clock = "none";
defparam \Mult0~mac .by_use_scan_in = "false";
defparam \Mult0~mac .bz_clock = "none";
defparam \Mult0~mac .coef_a_0 = 0;
defparam \Mult0~mac .coef_a_1 = 0;
defparam \Mult0~mac .coef_a_2 = 0;
defparam \Mult0~mac .coef_a_3 = 0;
defparam \Mult0~mac .coef_a_4 = 0;
defparam \Mult0~mac .coef_a_5 = 0;
defparam \Mult0~mac .coef_a_6 = 0;
defparam \Mult0~mac .coef_a_7 = 0;
defparam \Mult0~mac .coef_b_0 = 0;
defparam \Mult0~mac .coef_b_1 = 0;
defparam \Mult0~mac .coef_b_2 = 0;
defparam \Mult0~mac .coef_b_3 = 0;
defparam \Mult0~mac .coef_b_4 = 0;
defparam \Mult0~mac .coef_b_5 = 0;
defparam \Mult0~mac .coef_b_6 = 0;
defparam \Mult0~mac .coef_b_7 = 0;
defparam \Mult0~mac .coef_sel_a_clock = "none";
defparam \Mult0~mac .coef_sel_b_clock = "none";
defparam \Mult0~mac .delay_scan_out_ay = "false";
defparam \Mult0~mac .delay_scan_out_by = "false";
defparam \Mult0~mac .enable_double_accum = "false";
defparam \Mult0~mac .load_const_clock = "none";
defparam \Mult0~mac .load_const_value = 0;
defparam \Mult0~mac .mode_sub_location = 0;
defparam \Mult0~mac .negate_clock = "none";
defparam \Mult0~mac .operand_source_max = "input";
defparam \Mult0~mac .operand_source_may = "input";
defparam \Mult0~mac .operand_source_mbx = "input";
defparam \Mult0~mac .operand_source_mby = "input";
defparam \Mult0~mac .operation_mode = "m18x18_full";
defparam \Mult0~mac .output_clock = "none";
defparam \Mult0~mac .preadder_subtract_a = "false";
defparam \Mult0~mac .preadder_subtract_b = "false";
defparam \Mult0~mac .result_a_width = 64;
defparam \Mult0~mac .signed_max = "false";
defparam \Mult0~mac .signed_may = "false";
defparam \Mult0~mac .signed_mbx = "false";
defparam \Mult0~mac .signed_mby = "false";
defparam \Mult0~mac .sub_clock = "none";
defparam \Mult0~mac .use_chainadder = "false";

endmodule

module first_nios2_system_ama_register_function_31 (
	data_in,
	aclr,
	ena,
	data_out_wire_6,
	data_out_wire_7,
	data_out_wire_8,
	data_out_wire_9,
	data_out_wire_15,
	data_out_wire_5,
	data_out_wire_12,
	data_out_wire_11,
	data_out_wire_10,
	data_out_wire_4,
	data_out_wire_3,
	data_out_wire_1,
	data_out_wire_14,
	data_out_wire_2,
	data_out_wire_0,
	data_out_wire_13,
	clock)/* synthesis synthesis_greybox=1 */;
input 	[33:0] data_in;
input 	[3:0] aclr;
input 	[3:0] ena;
output 	data_out_wire_6;
output 	data_out_wire_7;
output 	data_out_wire_8;
output 	data_out_wire_9;
output 	data_out_wire_15;
output 	data_out_wire_5;
output 	data_out_wire_12;
output 	data_out_wire_11;
output 	data_out_wire_10;
output 	data_out_wire_4;
output 	data_out_wire_3;
output 	data_out_wire_1;
output 	data_out_wire_14;
output 	data_out_wire_2;
output 	data_out_wire_0;
output 	data_out_wire_13;
input 	[3:0] clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \data_out_wire[6] (
	.clk(clock[0]),
	.d(data_in[6]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!ena[0]),
	.q(data_out_wire_6),
	.prn(vcc));
defparam \data_out_wire[6] .is_wysiwyg = "true";
defparam \data_out_wire[6] .power_up = "low";

dffeas \data_out_wire[7] (
	.clk(clock[0]),
	.d(data_in[7]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!ena[0]),
	.q(data_out_wire_7),
	.prn(vcc));
defparam \data_out_wire[7] .is_wysiwyg = "true";
defparam \data_out_wire[7] .power_up = "low";

dffeas \data_out_wire[8] (
	.clk(clock[0]),
	.d(data_in[8]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!ena[0]),
	.q(data_out_wire_8),
	.prn(vcc));
defparam \data_out_wire[8] .is_wysiwyg = "true";
defparam \data_out_wire[8] .power_up = "low";

dffeas \data_out_wire[9] (
	.clk(clock[0]),
	.d(data_in[9]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!ena[0]),
	.q(data_out_wire_9),
	.prn(vcc));
defparam \data_out_wire[9] .is_wysiwyg = "true";
defparam \data_out_wire[9] .power_up = "low";

dffeas \data_out_wire[15] (
	.clk(clock[0]),
	.d(data_in[15]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!ena[0]),
	.q(data_out_wire_15),
	.prn(vcc));
defparam \data_out_wire[15] .is_wysiwyg = "true";
defparam \data_out_wire[15] .power_up = "low";

dffeas \data_out_wire[5] (
	.clk(clock[0]),
	.d(data_in[5]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!ena[0]),
	.q(data_out_wire_5),
	.prn(vcc));
defparam \data_out_wire[5] .is_wysiwyg = "true";
defparam \data_out_wire[5] .power_up = "low";

dffeas \data_out_wire[12] (
	.clk(clock[0]),
	.d(data_in[12]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!ena[0]),
	.q(data_out_wire_12),
	.prn(vcc));
defparam \data_out_wire[12] .is_wysiwyg = "true";
defparam \data_out_wire[12] .power_up = "low";

dffeas \data_out_wire[11] (
	.clk(clock[0]),
	.d(data_in[11]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!ena[0]),
	.q(data_out_wire_11),
	.prn(vcc));
defparam \data_out_wire[11] .is_wysiwyg = "true";
defparam \data_out_wire[11] .power_up = "low";

dffeas \data_out_wire[10] (
	.clk(clock[0]),
	.d(data_in[10]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!ena[0]),
	.q(data_out_wire_10),
	.prn(vcc));
defparam \data_out_wire[10] .is_wysiwyg = "true";
defparam \data_out_wire[10] .power_up = "low";

dffeas \data_out_wire[4] (
	.clk(clock[0]),
	.d(data_in[4]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!ena[0]),
	.q(data_out_wire_4),
	.prn(vcc));
defparam \data_out_wire[4] .is_wysiwyg = "true";
defparam \data_out_wire[4] .power_up = "low";

dffeas \data_out_wire[3] (
	.clk(clock[0]),
	.d(data_in[3]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!ena[0]),
	.q(data_out_wire_3),
	.prn(vcc));
defparam \data_out_wire[3] .is_wysiwyg = "true";
defparam \data_out_wire[3] .power_up = "low";

dffeas \data_out_wire[1] (
	.clk(clock[0]),
	.d(data_in[1]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!ena[0]),
	.q(data_out_wire_1),
	.prn(vcc));
defparam \data_out_wire[1] .is_wysiwyg = "true";
defparam \data_out_wire[1] .power_up = "low";

dffeas \data_out_wire[14] (
	.clk(clock[0]),
	.d(data_in[14]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!ena[0]),
	.q(data_out_wire_14),
	.prn(vcc));
defparam \data_out_wire[14] .is_wysiwyg = "true";
defparam \data_out_wire[14] .power_up = "low";

dffeas \data_out_wire[2] (
	.clk(clock[0]),
	.d(data_in[2]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!ena[0]),
	.q(data_out_wire_2),
	.prn(vcc));
defparam \data_out_wire[2] .is_wysiwyg = "true";
defparam \data_out_wire[2] .power_up = "low";

dffeas \data_out_wire[0] (
	.clk(clock[0]),
	.d(data_in[0]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!ena[0]),
	.q(data_out_wire_0),
	.prn(vcc));
defparam \data_out_wire[0] .is_wysiwyg = "true";
defparam \data_out_wire[0] .power_up = "low";

dffeas \data_out_wire[13] (
	.clk(clock[0]),
	.d(data_in[13]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!ena[0]),
	.q(data_out_wire_13),
	.prn(vcc));
defparam \data_out_wire[13] .is_wysiwyg = "true";
defparam \data_out_wire[13] .power_up = "low";

endmodule

module first_nios2_system_altera_mult_add_2 (
	E_src1_22,
	E_src1_23,
	E_src1_24,
	E_src1_25,
	E_src1_31,
	E_src2_7,
	E_src1_21,
	E_src2_11,
	E_src1_28,
	E_src2_10,
	E_src1_27,
	E_src2_8,
	E_src2_9,
	E_src2_5,
	E_src2_6,
	E_src1_26,
	E_src1_20,
	E_src1_19,
	E_src1_17,
	E_src1_30,
	E_src1_18,
	E_src1_16,
	E_src2_15,
	E_src2_12,
	E_src2_13,
	E_src2_14,
	E_src1_29,
	r_sync_rst,
	A_mem_stall,
	E_src2_3,
	E_src2_0,
	E_src2_2,
	E_src2_4,
	E_src2_1,
	data_out_wire_6,
	data_out_wire_7,
	data_out_wire_8,
	data_out_wire_9,
	data_out_wire_15,
	data_out_wire_5,
	data_out_wire_12,
	data_out_wire_11,
	data_out_wire_10,
	data_out_wire_4,
	data_out_wire_3,
	data_out_wire_1,
	data_out_wire_14,
	data_out_wire_2,
	data_out_wire_0,
	data_out_wire_13,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	E_src1_22;
input 	E_src1_23;
input 	E_src1_24;
input 	E_src1_25;
input 	E_src1_31;
input 	E_src2_7;
input 	E_src1_21;
input 	E_src2_11;
input 	E_src1_28;
input 	E_src2_10;
input 	E_src1_27;
input 	E_src2_8;
input 	E_src2_9;
input 	E_src2_5;
input 	E_src2_6;
input 	E_src1_26;
input 	E_src1_20;
input 	E_src1_19;
input 	E_src1_17;
input 	E_src1_30;
input 	E_src1_18;
input 	E_src1_16;
input 	E_src2_15;
input 	E_src2_12;
input 	E_src2_13;
input 	E_src2_14;
input 	E_src1_29;
input 	r_sync_rst;
input 	A_mem_stall;
input 	E_src2_3;
input 	E_src2_0;
input 	E_src2_2;
input 	E_src2_4;
input 	E_src2_1;
output 	data_out_wire_6;
output 	data_out_wire_7;
output 	data_out_wire_8;
output 	data_out_wire_9;
output 	data_out_wire_15;
output 	data_out_wire_5;
output 	data_out_wire_12;
output 	data_out_wire_11;
output 	data_out_wire_10;
output 	data_out_wire_4;
output 	data_out_wire_3;
output 	data_out_wire_1;
output 	data_out_wire_14;
output 	data_out_wire_2;
output 	data_out_wire_0;
output 	data_out_wire_13;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



first_nios2_system_altera_mult_add_37p2_2 auto_generated(
	.E_src1_22(E_src1_22),
	.E_src1_23(E_src1_23),
	.E_src1_24(E_src1_24),
	.E_src1_25(E_src1_25),
	.E_src1_31(E_src1_31),
	.E_src2_7(E_src2_7),
	.E_src1_21(E_src1_21),
	.E_src2_11(E_src2_11),
	.E_src1_28(E_src1_28),
	.E_src2_10(E_src2_10),
	.E_src1_27(E_src1_27),
	.E_src2_8(E_src2_8),
	.E_src2_9(E_src2_9),
	.E_src2_5(E_src2_5),
	.E_src2_6(E_src2_6),
	.E_src1_26(E_src1_26),
	.E_src1_20(E_src1_20),
	.E_src1_19(E_src1_19),
	.E_src1_17(E_src1_17),
	.E_src1_30(E_src1_30),
	.E_src1_18(E_src1_18),
	.E_src1_16(E_src1_16),
	.E_src2_15(E_src2_15),
	.E_src2_12(E_src2_12),
	.E_src2_13(E_src2_13),
	.E_src2_14(E_src2_14),
	.E_src1_29(E_src1_29),
	.r_sync_rst(r_sync_rst),
	.A_mem_stall(A_mem_stall),
	.E_src2_3(E_src2_3),
	.E_src2_0(E_src2_0),
	.E_src2_2(E_src2_2),
	.E_src2_4(E_src2_4),
	.E_src2_1(E_src2_1),
	.data_out_wire_6(data_out_wire_6),
	.data_out_wire_7(data_out_wire_7),
	.data_out_wire_8(data_out_wire_8),
	.data_out_wire_9(data_out_wire_9),
	.data_out_wire_15(data_out_wire_15),
	.data_out_wire_5(data_out_wire_5),
	.data_out_wire_12(data_out_wire_12),
	.data_out_wire_11(data_out_wire_11),
	.data_out_wire_10(data_out_wire_10),
	.data_out_wire_4(data_out_wire_4),
	.data_out_wire_3(data_out_wire_3),
	.data_out_wire_1(data_out_wire_1),
	.data_out_wire_14(data_out_wire_14),
	.data_out_wire_2(data_out_wire_2),
	.data_out_wire_0(data_out_wire_0),
	.data_out_wire_13(data_out_wire_13),
	.clk_clk(clk_clk));

endmodule

module first_nios2_system_altera_mult_add_37p2_2 (
	E_src1_22,
	E_src1_23,
	E_src1_24,
	E_src1_25,
	E_src1_31,
	E_src2_7,
	E_src1_21,
	E_src2_11,
	E_src1_28,
	E_src2_10,
	E_src1_27,
	E_src2_8,
	E_src2_9,
	E_src2_5,
	E_src2_6,
	E_src1_26,
	E_src1_20,
	E_src1_19,
	E_src1_17,
	E_src1_30,
	E_src1_18,
	E_src1_16,
	E_src2_15,
	E_src2_12,
	E_src2_13,
	E_src2_14,
	E_src1_29,
	r_sync_rst,
	A_mem_stall,
	E_src2_3,
	E_src2_0,
	E_src2_2,
	E_src2_4,
	E_src2_1,
	data_out_wire_6,
	data_out_wire_7,
	data_out_wire_8,
	data_out_wire_9,
	data_out_wire_15,
	data_out_wire_5,
	data_out_wire_12,
	data_out_wire_11,
	data_out_wire_10,
	data_out_wire_4,
	data_out_wire_3,
	data_out_wire_1,
	data_out_wire_14,
	data_out_wire_2,
	data_out_wire_0,
	data_out_wire_13,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	E_src1_22;
input 	E_src1_23;
input 	E_src1_24;
input 	E_src1_25;
input 	E_src1_31;
input 	E_src2_7;
input 	E_src1_21;
input 	E_src2_11;
input 	E_src1_28;
input 	E_src2_10;
input 	E_src1_27;
input 	E_src2_8;
input 	E_src2_9;
input 	E_src2_5;
input 	E_src2_6;
input 	E_src1_26;
input 	E_src1_20;
input 	E_src1_19;
input 	E_src1_17;
input 	E_src1_30;
input 	E_src1_18;
input 	E_src1_16;
input 	E_src2_15;
input 	E_src2_12;
input 	E_src2_13;
input 	E_src2_14;
input 	E_src1_29;
input 	r_sync_rst;
input 	A_mem_stall;
input 	E_src2_3;
input 	E_src2_0;
input 	E_src2_2;
input 	E_src2_4;
input 	E_src2_1;
output 	data_out_wire_6;
output 	data_out_wire_7;
output 	data_out_wire_8;
output 	data_out_wire_9;
output 	data_out_wire_15;
output 	data_out_wire_5;
output 	data_out_wire_12;
output 	data_out_wire_11;
output 	data_out_wire_10;
output 	data_out_wire_4;
output 	data_out_wire_3;
output 	data_out_wire_1;
output 	data_out_wire_14;
output 	data_out_wire_2;
output 	data_out_wire_0;
output 	data_out_wire_13;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



first_nios2_system_altera_mult_add_rtl_3 altera_mult_add_rtl1(
	.E_src1_22(E_src1_22),
	.E_src1_23(E_src1_23),
	.E_src1_24(E_src1_24),
	.E_src1_25(E_src1_25),
	.E_src1_31(E_src1_31),
	.E_src2_7(E_src2_7),
	.E_src1_21(E_src1_21),
	.E_src2_11(E_src2_11),
	.E_src1_28(E_src1_28),
	.E_src2_10(E_src2_10),
	.E_src1_27(E_src1_27),
	.E_src2_8(E_src2_8),
	.E_src2_9(E_src2_9),
	.E_src2_5(E_src2_5),
	.E_src2_6(E_src2_6),
	.E_src1_26(E_src1_26),
	.E_src1_20(E_src1_20),
	.E_src1_19(E_src1_19),
	.E_src1_17(E_src1_17),
	.E_src1_30(E_src1_30),
	.E_src1_18(E_src1_18),
	.E_src1_16(E_src1_16),
	.E_src2_15(E_src2_15),
	.E_src2_12(E_src2_12),
	.E_src2_13(E_src2_13),
	.E_src2_14(E_src2_14),
	.E_src1_29(E_src1_29),
	.r_sync_rst(r_sync_rst),
	.A_mem_stall(A_mem_stall),
	.E_src2_3(E_src2_3),
	.E_src2_0(E_src2_0),
	.E_src2_2(E_src2_2),
	.E_src2_4(E_src2_4),
	.E_src2_1(E_src2_1),
	.data_out_wire_6(data_out_wire_6),
	.data_out_wire_7(data_out_wire_7),
	.data_out_wire_8(data_out_wire_8),
	.data_out_wire_9(data_out_wire_9),
	.data_out_wire_15(data_out_wire_15),
	.data_out_wire_5(data_out_wire_5),
	.data_out_wire_12(data_out_wire_12),
	.data_out_wire_11(data_out_wire_11),
	.data_out_wire_10(data_out_wire_10),
	.data_out_wire_4(data_out_wire_4),
	.data_out_wire_3(data_out_wire_3),
	.data_out_wire_1(data_out_wire_1),
	.data_out_wire_14(data_out_wire_14),
	.data_out_wire_2(data_out_wire_2),
	.data_out_wire_0(data_out_wire_0),
	.data_out_wire_13(data_out_wire_13),
	.clk_clk(clk_clk));

endmodule

module first_nios2_system_altera_mult_add_rtl_3 (
	E_src1_22,
	E_src1_23,
	E_src1_24,
	E_src1_25,
	E_src1_31,
	E_src2_7,
	E_src1_21,
	E_src2_11,
	E_src1_28,
	E_src2_10,
	E_src1_27,
	E_src2_8,
	E_src2_9,
	E_src2_5,
	E_src2_6,
	E_src1_26,
	E_src1_20,
	E_src1_19,
	E_src1_17,
	E_src1_30,
	E_src1_18,
	E_src1_16,
	E_src2_15,
	E_src2_12,
	E_src2_13,
	E_src2_14,
	E_src1_29,
	r_sync_rst,
	A_mem_stall,
	E_src2_3,
	E_src2_0,
	E_src2_2,
	E_src2_4,
	E_src2_1,
	data_out_wire_6,
	data_out_wire_7,
	data_out_wire_8,
	data_out_wire_9,
	data_out_wire_15,
	data_out_wire_5,
	data_out_wire_12,
	data_out_wire_11,
	data_out_wire_10,
	data_out_wire_4,
	data_out_wire_3,
	data_out_wire_1,
	data_out_wire_14,
	data_out_wire_2,
	data_out_wire_0,
	data_out_wire_13,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	E_src1_22;
input 	E_src1_23;
input 	E_src1_24;
input 	E_src1_25;
input 	E_src1_31;
input 	E_src2_7;
input 	E_src1_21;
input 	E_src2_11;
input 	E_src1_28;
input 	E_src2_10;
input 	E_src1_27;
input 	E_src2_8;
input 	E_src2_9;
input 	E_src2_5;
input 	E_src2_6;
input 	E_src1_26;
input 	E_src1_20;
input 	E_src1_19;
input 	E_src1_17;
input 	E_src1_30;
input 	E_src1_18;
input 	E_src1_16;
input 	E_src2_15;
input 	E_src2_12;
input 	E_src2_13;
input 	E_src2_14;
input 	E_src1_29;
input 	r_sync_rst;
input 	A_mem_stall;
input 	E_src2_3;
input 	E_src2_0;
input 	E_src2_2;
input 	E_src2_4;
input 	E_src2_1;
output 	data_out_wire_6;
output 	data_out_wire_7;
output 	data_out_wire_8;
output 	data_out_wire_9;
output 	data_out_wire_15;
output 	data_out_wire_5;
output 	data_out_wire_12;
output 	data_out_wire_11;
output 	data_out_wire_10;
output 	data_out_wire_4;
output 	data_out_wire_3;
output 	data_out_wire_1;
output 	data_out_wire_14;
output 	data_out_wire_2;
output 	data_out_wire_0;
output 	data_out_wire_13;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



first_nios2_system_ama_multiplier_function_2 multiplier_block(
	.E_src1_22(E_src1_22),
	.E_src1_23(E_src1_23),
	.E_src1_24(E_src1_24),
	.E_src1_25(E_src1_25),
	.E_src1_31(E_src1_31),
	.E_src2_7(E_src2_7),
	.E_src1_21(E_src1_21),
	.E_src2_11(E_src2_11),
	.E_src1_28(E_src1_28),
	.E_src2_10(E_src2_10),
	.E_src1_27(E_src1_27),
	.E_src2_8(E_src2_8),
	.E_src2_9(E_src2_9),
	.E_src2_5(E_src2_5),
	.E_src2_6(E_src2_6),
	.E_src1_26(E_src1_26),
	.E_src1_20(E_src1_20),
	.E_src1_19(E_src1_19),
	.E_src1_17(E_src1_17),
	.E_src1_30(E_src1_30),
	.E_src1_18(E_src1_18),
	.E_src1_16(E_src1_16),
	.E_src2_15(E_src2_15),
	.E_src2_12(E_src2_12),
	.E_src2_13(E_src2_13),
	.E_src2_14(E_src2_14),
	.E_src1_29(E_src1_29),
	.r_sync_rst(r_sync_rst),
	.A_mem_stall(A_mem_stall),
	.E_src2_3(E_src2_3),
	.E_src2_0(E_src2_0),
	.E_src2_2(E_src2_2),
	.E_src2_4(E_src2_4),
	.E_src2_1(E_src2_1),
	.data_out_wire_6(data_out_wire_6),
	.data_out_wire_7(data_out_wire_7),
	.data_out_wire_8(data_out_wire_8),
	.data_out_wire_9(data_out_wire_9),
	.data_out_wire_15(data_out_wire_15),
	.data_out_wire_5(data_out_wire_5),
	.data_out_wire_12(data_out_wire_12),
	.data_out_wire_11(data_out_wire_11),
	.data_out_wire_10(data_out_wire_10),
	.data_out_wire_4(data_out_wire_4),
	.data_out_wire_3(data_out_wire_3),
	.data_out_wire_1(data_out_wire_1),
	.data_out_wire_14(data_out_wire_14),
	.data_out_wire_2(data_out_wire_2),
	.data_out_wire_0(data_out_wire_0),
	.data_out_wire_13(data_out_wire_13),
	.clk_clk(clk_clk));

endmodule

module first_nios2_system_ama_multiplier_function_2 (
	E_src1_22,
	E_src1_23,
	E_src1_24,
	E_src1_25,
	E_src1_31,
	E_src2_7,
	E_src1_21,
	E_src2_11,
	E_src1_28,
	E_src2_10,
	E_src1_27,
	E_src2_8,
	E_src2_9,
	E_src2_5,
	E_src2_6,
	E_src1_26,
	E_src1_20,
	E_src1_19,
	E_src1_17,
	E_src1_30,
	E_src1_18,
	E_src1_16,
	E_src2_15,
	E_src2_12,
	E_src2_13,
	E_src2_14,
	E_src1_29,
	r_sync_rst,
	A_mem_stall,
	E_src2_3,
	E_src2_0,
	E_src2_2,
	E_src2_4,
	E_src2_1,
	data_out_wire_6,
	data_out_wire_7,
	data_out_wire_8,
	data_out_wire_9,
	data_out_wire_15,
	data_out_wire_5,
	data_out_wire_12,
	data_out_wire_11,
	data_out_wire_10,
	data_out_wire_4,
	data_out_wire_3,
	data_out_wire_1,
	data_out_wire_14,
	data_out_wire_2,
	data_out_wire_0,
	data_out_wire_13,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	E_src1_22;
input 	E_src1_23;
input 	E_src1_24;
input 	E_src1_25;
input 	E_src1_31;
input 	E_src2_7;
input 	E_src1_21;
input 	E_src2_11;
input 	E_src1_28;
input 	E_src2_10;
input 	E_src1_27;
input 	E_src2_8;
input 	E_src2_9;
input 	E_src2_5;
input 	E_src2_6;
input 	E_src1_26;
input 	E_src1_20;
input 	E_src1_19;
input 	E_src1_17;
input 	E_src1_30;
input 	E_src1_18;
input 	E_src1_16;
input 	E_src2_15;
input 	E_src2_12;
input 	E_src2_13;
input 	E_src2_14;
input 	E_src1_29;
input 	r_sync_rst;
input 	A_mem_stall;
input 	E_src2_3;
input 	E_src2_0;
input 	E_src2_2;
input 	E_src2_4;
input 	E_src2_1;
output 	data_out_wire_6;
output 	data_out_wire_7;
output 	data_out_wire_8;
output 	data_out_wire_9;
output 	data_out_wire_15;
output 	data_out_wire_5;
output 	data_out_wire_12;
output 	data_out_wire_11;
output 	data_out_wire_10;
output 	data_out_wire_4;
output 	data_out_wire_3;
output 	data_out_wire_1;
output 	data_out_wire_14;
output 	data_out_wire_2;
output 	data_out_wire_0;
output 	data_out_wire_13;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \data_out_wire_0[0] ;
wire \data_out_wire_0[1] ;
wire \data_out_wire_0[2] ;
wire \data_out_wire_0[3] ;
wire \data_out_wire_0[4] ;
wire \data_out_wire_0[5] ;
wire \data_out_wire_0[6] ;
wire \data_out_wire_0[7] ;
wire \data_out_wire_0[8] ;
wire \data_out_wire_0[9] ;
wire \data_out_wire_0[10] ;
wire \data_out_wire_0[11] ;
wire \data_out_wire_0[12] ;
wire \data_out_wire_0[13] ;
wire \data_out_wire_0[14] ;
wire \data_out_wire_0[15] ;
wire \Mult0~8 ;
wire \Mult0~9 ;
wire \Mult0~10 ;
wire \Mult0~11 ;
wire \Mult0~12 ;
wire \Mult0~13 ;
wire \Mult0~14 ;
wire \Mult0~15 ;
wire \Mult0~16 ;
wire \Mult0~17 ;
wire \Mult0~18 ;
wire \Mult0~19 ;
wire \Mult0~20 ;
wire \Mult0~21 ;
wire \Mult0~22 ;
wire \Mult0~23 ;
wire \Mult0~24 ;
wire \Mult0~25 ;
wire \Mult0~26 ;
wire \Mult0~27 ;
wire \Mult0~28 ;
wire \Mult0~29 ;
wire \Mult0~30 ;
wire \Mult0~31 ;
wire \Mult0~32 ;
wire \Mult0~33 ;
wire \Mult0~34 ;
wire \Mult0~35 ;
wire \Mult0~36 ;
wire \Mult0~37 ;
wire \Mult0~38 ;
wire \Mult0~39 ;
wire \Mult0~40 ;
wire \Mult0~41 ;
wire \Mult0~42 ;
wire \Mult0~43 ;
wire \Mult0~44 ;
wire \Mult0~45 ;
wire \Mult0~46 ;
wire \Mult0~47 ;
wire \Mult0~48 ;
wire \Mult0~49 ;
wire \Mult0~50 ;
wire \Mult0~51 ;
wire \Mult0~52 ;
wire \Mult0~53 ;
wire \Mult0~54 ;
wire \Mult0~55 ;

wire [63:0] \Mult0~mac_RESULTA_bus ;

assign \data_out_wire_0[0]  = \Mult0~mac_RESULTA_bus [0];
assign \data_out_wire_0[1]  = \Mult0~mac_RESULTA_bus [1];
assign \data_out_wire_0[2]  = \Mult0~mac_RESULTA_bus [2];
assign \data_out_wire_0[3]  = \Mult0~mac_RESULTA_bus [3];
assign \data_out_wire_0[4]  = \Mult0~mac_RESULTA_bus [4];
assign \data_out_wire_0[5]  = \Mult0~mac_RESULTA_bus [5];
assign \data_out_wire_0[6]  = \Mult0~mac_RESULTA_bus [6];
assign \data_out_wire_0[7]  = \Mult0~mac_RESULTA_bus [7];
assign \data_out_wire_0[8]  = \Mult0~mac_RESULTA_bus [8];
assign \data_out_wire_0[9]  = \Mult0~mac_RESULTA_bus [9];
assign \data_out_wire_0[10]  = \Mult0~mac_RESULTA_bus [10];
assign \data_out_wire_0[11]  = \Mult0~mac_RESULTA_bus [11];
assign \data_out_wire_0[12]  = \Mult0~mac_RESULTA_bus [12];
assign \data_out_wire_0[13]  = \Mult0~mac_RESULTA_bus [13];
assign \data_out_wire_0[14]  = \Mult0~mac_RESULTA_bus [14];
assign \data_out_wire_0[15]  = \Mult0~mac_RESULTA_bus [15];
assign \Mult0~8  = \Mult0~mac_RESULTA_bus [16];
assign \Mult0~9  = \Mult0~mac_RESULTA_bus [17];
assign \Mult0~10  = \Mult0~mac_RESULTA_bus [18];
assign \Mult0~11  = \Mult0~mac_RESULTA_bus [19];
assign \Mult0~12  = \Mult0~mac_RESULTA_bus [20];
assign \Mult0~13  = \Mult0~mac_RESULTA_bus [21];
assign \Mult0~14  = \Mult0~mac_RESULTA_bus [22];
assign \Mult0~15  = \Mult0~mac_RESULTA_bus [23];
assign \Mult0~16  = \Mult0~mac_RESULTA_bus [24];
assign \Mult0~17  = \Mult0~mac_RESULTA_bus [25];
assign \Mult0~18  = \Mult0~mac_RESULTA_bus [26];
assign \Mult0~19  = \Mult0~mac_RESULTA_bus [27];
assign \Mult0~20  = \Mult0~mac_RESULTA_bus [28];
assign \Mult0~21  = \Mult0~mac_RESULTA_bus [29];
assign \Mult0~22  = \Mult0~mac_RESULTA_bus [30];
assign \Mult0~23  = \Mult0~mac_RESULTA_bus [31];
assign \Mult0~24  = \Mult0~mac_RESULTA_bus [32];
assign \Mult0~25  = \Mult0~mac_RESULTA_bus [33];
assign \Mult0~26  = \Mult0~mac_RESULTA_bus [34];
assign \Mult0~27  = \Mult0~mac_RESULTA_bus [35];
assign \Mult0~28  = \Mult0~mac_RESULTA_bus [36];
assign \Mult0~29  = \Mult0~mac_RESULTA_bus [37];
assign \Mult0~30  = \Mult0~mac_RESULTA_bus [38];
assign \Mult0~31  = \Mult0~mac_RESULTA_bus [39];
assign \Mult0~32  = \Mult0~mac_RESULTA_bus [40];
assign \Mult0~33  = \Mult0~mac_RESULTA_bus [41];
assign \Mult0~34  = \Mult0~mac_RESULTA_bus [42];
assign \Mult0~35  = \Mult0~mac_RESULTA_bus [43];
assign \Mult0~36  = \Mult0~mac_RESULTA_bus [44];
assign \Mult0~37  = \Mult0~mac_RESULTA_bus [45];
assign \Mult0~38  = \Mult0~mac_RESULTA_bus [46];
assign \Mult0~39  = \Mult0~mac_RESULTA_bus [47];
assign \Mult0~40  = \Mult0~mac_RESULTA_bus [48];
assign \Mult0~41  = \Mult0~mac_RESULTA_bus [49];
assign \Mult0~42  = \Mult0~mac_RESULTA_bus [50];
assign \Mult0~43  = \Mult0~mac_RESULTA_bus [51];
assign \Mult0~44  = \Mult0~mac_RESULTA_bus [52];
assign \Mult0~45  = \Mult0~mac_RESULTA_bus [53];
assign \Mult0~46  = \Mult0~mac_RESULTA_bus [54];
assign \Mult0~47  = \Mult0~mac_RESULTA_bus [55];
assign \Mult0~48  = \Mult0~mac_RESULTA_bus [56];
assign \Mult0~49  = \Mult0~mac_RESULTA_bus [57];
assign \Mult0~50  = \Mult0~mac_RESULTA_bus [58];
assign \Mult0~51  = \Mult0~mac_RESULTA_bus [59];
assign \Mult0~52  = \Mult0~mac_RESULTA_bus [60];
assign \Mult0~53  = \Mult0~mac_RESULTA_bus [61];
assign \Mult0~54  = \Mult0~mac_RESULTA_bus [62];
assign \Mult0~55  = \Mult0~mac_RESULTA_bus [63];

first_nios2_system_ama_register_function_50 multiplier_register_block_0(
	.data_in({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\data_out_wire_0[15] ,\data_out_wire_0[14] ,\data_out_wire_0[13] ,\data_out_wire_0[12] ,\data_out_wire_0[11] ,\data_out_wire_0[10] ,\data_out_wire_0[9] ,\data_out_wire_0[8] ,\data_out_wire_0[7] ,
\data_out_wire_0[6] ,\data_out_wire_0[5] ,\data_out_wire_0[4] ,\data_out_wire_0[3] ,\data_out_wire_0[2] ,\data_out_wire_0[1] ,\data_out_wire_0[0] }),
	.aclr({gnd,gnd,gnd,r_sync_rst}),
	.ena({gnd,gnd,gnd,A_mem_stall}),
	.data_out_wire_6(data_out_wire_6),
	.data_out_wire_7(data_out_wire_7),
	.data_out_wire_8(data_out_wire_8),
	.data_out_wire_9(data_out_wire_9),
	.data_out_wire_15(data_out_wire_15),
	.data_out_wire_5(data_out_wire_5),
	.data_out_wire_12(data_out_wire_12),
	.data_out_wire_11(data_out_wire_11),
	.data_out_wire_10(data_out_wire_10),
	.data_out_wire_4(data_out_wire_4),
	.data_out_wire_3(data_out_wire_3),
	.data_out_wire_1(data_out_wire_1),
	.data_out_wire_14(data_out_wire_14),
	.data_out_wire_2(data_out_wire_2),
	.data_out_wire_0(data_out_wire_0),
	.data_out_wire_13(data_out_wire_13),
	.clock({gnd,gnd,gnd,clk_clk}));

cyclonev_mac \Mult0~mac (
	.sub(gnd),
	.negate(gnd),
	.accumulate(gnd),
	.loadconst(gnd),
	.ax({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,E_src2_15,E_src2_14,E_src2_13,E_src2_12,E_src2_11,E_src2_10,E_src2_9,E_src2_8,E_src2_7,E_src2_6,E_src2_5,E_src2_4,E_src2_3,E_src2_2,E_src2_1,E_src2_0}),
	.ay({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,E_src1_31,E_src1_30,E_src1_29,E_src1_28,E_src1_27,E_src1_26,E_src1_25,E_src1_24,E_src1_23,E_src1_22,E_src1_21,E_src1_20,E_src1_19,E_src1_18,E_src1_17,E_src1_16}),
	.az(26'b00000000000000000000000000),
	.bx(18'b000000000000000000),
	.by(19'b0000000000000000000),
	.bz(18'b000000000000000000),
	.coefsela(3'b000),
	.coefselb(3'b000),
	.clk(3'b000),
	.aclr(2'b00),
	.ena(3'b111),
	.scanin(27'b000000000000000000000000000),
	.chainin(1'b0),
	.dftout(),
	.resulta(\Mult0~mac_RESULTA_bus ),
	.resultb(),
	.scanout(),
	.chainout());
defparam \Mult0~mac .accumulate_clock = "none";
defparam \Mult0~mac .ax_clock = "none";
defparam \Mult0~mac .ax_width = 16;
defparam \Mult0~mac .ay_scan_in_clock = "none";
defparam \Mult0~mac .ay_scan_in_width = 16;
defparam \Mult0~mac .ay_use_scan_in = "false";
defparam \Mult0~mac .az_clock = "none";
defparam \Mult0~mac .bx_clock = "none";
defparam \Mult0~mac .by_clock = "none";
defparam \Mult0~mac .by_use_scan_in = "false";
defparam \Mult0~mac .bz_clock = "none";
defparam \Mult0~mac .coef_a_0 = 0;
defparam \Mult0~mac .coef_a_1 = 0;
defparam \Mult0~mac .coef_a_2 = 0;
defparam \Mult0~mac .coef_a_3 = 0;
defparam \Mult0~mac .coef_a_4 = 0;
defparam \Mult0~mac .coef_a_5 = 0;
defparam \Mult0~mac .coef_a_6 = 0;
defparam \Mult0~mac .coef_a_7 = 0;
defparam \Mult0~mac .coef_b_0 = 0;
defparam \Mult0~mac .coef_b_1 = 0;
defparam \Mult0~mac .coef_b_2 = 0;
defparam \Mult0~mac .coef_b_3 = 0;
defparam \Mult0~mac .coef_b_4 = 0;
defparam \Mult0~mac .coef_b_5 = 0;
defparam \Mult0~mac .coef_b_6 = 0;
defparam \Mult0~mac .coef_b_7 = 0;
defparam \Mult0~mac .coef_sel_a_clock = "none";
defparam \Mult0~mac .coef_sel_b_clock = "none";
defparam \Mult0~mac .delay_scan_out_ay = "false";
defparam \Mult0~mac .delay_scan_out_by = "false";
defparam \Mult0~mac .enable_double_accum = "false";
defparam \Mult0~mac .load_const_clock = "none";
defparam \Mult0~mac .load_const_value = 0;
defparam \Mult0~mac .mode_sub_location = 0;
defparam \Mult0~mac .negate_clock = "none";
defparam \Mult0~mac .operand_source_max = "input";
defparam \Mult0~mac .operand_source_may = "input";
defparam \Mult0~mac .operand_source_mbx = "input";
defparam \Mult0~mac .operand_source_mby = "input";
defparam \Mult0~mac .operation_mode = "m18x18_full";
defparam \Mult0~mac .output_clock = "none";
defparam \Mult0~mac .preadder_subtract_a = "false";
defparam \Mult0~mac .preadder_subtract_b = "false";
defparam \Mult0~mac .result_a_width = 64;
defparam \Mult0~mac .signed_max = "false";
defparam \Mult0~mac .signed_may = "false";
defparam \Mult0~mac .signed_mbx = "false";
defparam \Mult0~mac .signed_mby = "false";
defparam \Mult0~mac .sub_clock = "none";
defparam \Mult0~mac .use_chainadder = "false";

endmodule

module first_nios2_system_ama_register_function_50 (
	data_in,
	aclr,
	ena,
	data_out_wire_6,
	data_out_wire_7,
	data_out_wire_8,
	data_out_wire_9,
	data_out_wire_15,
	data_out_wire_5,
	data_out_wire_12,
	data_out_wire_11,
	data_out_wire_10,
	data_out_wire_4,
	data_out_wire_3,
	data_out_wire_1,
	data_out_wire_14,
	data_out_wire_2,
	data_out_wire_0,
	data_out_wire_13,
	clock)/* synthesis synthesis_greybox=1 */;
input 	[33:0] data_in;
input 	[3:0] aclr;
input 	[3:0] ena;
output 	data_out_wire_6;
output 	data_out_wire_7;
output 	data_out_wire_8;
output 	data_out_wire_9;
output 	data_out_wire_15;
output 	data_out_wire_5;
output 	data_out_wire_12;
output 	data_out_wire_11;
output 	data_out_wire_10;
output 	data_out_wire_4;
output 	data_out_wire_3;
output 	data_out_wire_1;
output 	data_out_wire_14;
output 	data_out_wire_2;
output 	data_out_wire_0;
output 	data_out_wire_13;
input 	[3:0] clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \data_out_wire[6] (
	.clk(clock[0]),
	.d(data_in[6]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!ena[0]),
	.q(data_out_wire_6),
	.prn(vcc));
defparam \data_out_wire[6] .is_wysiwyg = "true";
defparam \data_out_wire[6] .power_up = "low";

dffeas \data_out_wire[7] (
	.clk(clock[0]),
	.d(data_in[7]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!ena[0]),
	.q(data_out_wire_7),
	.prn(vcc));
defparam \data_out_wire[7] .is_wysiwyg = "true";
defparam \data_out_wire[7] .power_up = "low";

dffeas \data_out_wire[8] (
	.clk(clock[0]),
	.d(data_in[8]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!ena[0]),
	.q(data_out_wire_8),
	.prn(vcc));
defparam \data_out_wire[8] .is_wysiwyg = "true";
defparam \data_out_wire[8] .power_up = "low";

dffeas \data_out_wire[9] (
	.clk(clock[0]),
	.d(data_in[9]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!ena[0]),
	.q(data_out_wire_9),
	.prn(vcc));
defparam \data_out_wire[9] .is_wysiwyg = "true";
defparam \data_out_wire[9] .power_up = "low";

dffeas \data_out_wire[15] (
	.clk(clock[0]),
	.d(data_in[15]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!ena[0]),
	.q(data_out_wire_15),
	.prn(vcc));
defparam \data_out_wire[15] .is_wysiwyg = "true";
defparam \data_out_wire[15] .power_up = "low";

dffeas \data_out_wire[5] (
	.clk(clock[0]),
	.d(data_in[5]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!ena[0]),
	.q(data_out_wire_5),
	.prn(vcc));
defparam \data_out_wire[5] .is_wysiwyg = "true";
defparam \data_out_wire[5] .power_up = "low";

dffeas \data_out_wire[12] (
	.clk(clock[0]),
	.d(data_in[12]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!ena[0]),
	.q(data_out_wire_12),
	.prn(vcc));
defparam \data_out_wire[12] .is_wysiwyg = "true";
defparam \data_out_wire[12] .power_up = "low";

dffeas \data_out_wire[11] (
	.clk(clock[0]),
	.d(data_in[11]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!ena[0]),
	.q(data_out_wire_11),
	.prn(vcc));
defparam \data_out_wire[11] .is_wysiwyg = "true";
defparam \data_out_wire[11] .power_up = "low";

dffeas \data_out_wire[10] (
	.clk(clock[0]),
	.d(data_in[10]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!ena[0]),
	.q(data_out_wire_10),
	.prn(vcc));
defparam \data_out_wire[10] .is_wysiwyg = "true";
defparam \data_out_wire[10] .power_up = "low";

dffeas \data_out_wire[4] (
	.clk(clock[0]),
	.d(data_in[4]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!ena[0]),
	.q(data_out_wire_4),
	.prn(vcc));
defparam \data_out_wire[4] .is_wysiwyg = "true";
defparam \data_out_wire[4] .power_up = "low";

dffeas \data_out_wire[3] (
	.clk(clock[0]),
	.d(data_in[3]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!ena[0]),
	.q(data_out_wire_3),
	.prn(vcc));
defparam \data_out_wire[3] .is_wysiwyg = "true";
defparam \data_out_wire[3] .power_up = "low";

dffeas \data_out_wire[1] (
	.clk(clock[0]),
	.d(data_in[1]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!ena[0]),
	.q(data_out_wire_1),
	.prn(vcc));
defparam \data_out_wire[1] .is_wysiwyg = "true";
defparam \data_out_wire[1] .power_up = "low";

dffeas \data_out_wire[14] (
	.clk(clock[0]),
	.d(data_in[14]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!ena[0]),
	.q(data_out_wire_14),
	.prn(vcc));
defparam \data_out_wire[14] .is_wysiwyg = "true";
defparam \data_out_wire[14] .power_up = "low";

dffeas \data_out_wire[2] (
	.clk(clock[0]),
	.d(data_in[2]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!ena[0]),
	.q(data_out_wire_2),
	.prn(vcc));
defparam \data_out_wire[2] .is_wysiwyg = "true";
defparam \data_out_wire[2] .power_up = "low";

dffeas \data_out_wire[0] (
	.clk(clock[0]),
	.d(data_in[0]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!ena[0]),
	.q(data_out_wire_0),
	.prn(vcc));
defparam \data_out_wire[0] .is_wysiwyg = "true";
defparam \data_out_wire[0] .power_up = "low";

dffeas \data_out_wire[13] (
	.clk(clock[0]),
	.d(data_in[13]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!ena[0]),
	.q(data_out_wire_13),
	.prn(vcc));
defparam \data_out_wire[13] .is_wysiwyg = "true";
defparam \data_out_wire[13] .power_up = "low";

endmodule

module first_nios2_system_first_nios2_system_cpu_cpu_nios2_oci (
	readdata_0,
	readdata_1,
	readdata_2,
	readdata_3,
	readdata_4,
	readdata_5,
	readdata_6,
	readdata_7,
	readdata_22,
	readdata_23,
	readdata_24,
	readdata_25,
	readdata_31,
	readdata_21,
	readdata_11,
	readdata_28,
	readdata_10,
	readdata_27,
	readdata_8,
	readdata_9,
	readdata_26,
	readdata_20,
	readdata_19,
	readdata_17,
	readdata_30,
	readdata_18,
	readdata_16,
	readdata_15,
	readdata_12,
	readdata_13,
	readdata_14,
	readdata_29,
	sr_0,
	ir_out_0,
	ir_out_1,
	d_write,
	r_sync_rst,
	W_debug_mode,
	oci_single_step_mode,
	jtag_break,
	saved_grant_0,
	waitrequest,
	mem_used_1,
	WideOr1,
	mem,
	oci_ienable_1,
	oci_ienable_16,
	writedata_nxt,
	address_nxt,
	debugaccess_nxt,
	r_early_rst,
	byteenable_nxt,
	altera_internal_jtag,
	altera_internal_jtag1,
	state_1,
	state_4,
	virtual_ir_scan_reg,
	state_3,
	state_8,
	splitter_nodes_receive_1_3,
	irf_reg_0_2,
	irf_reg_1_2,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	readdata_0;
output 	readdata_1;
output 	readdata_2;
output 	readdata_3;
output 	readdata_4;
output 	readdata_5;
output 	readdata_6;
output 	readdata_7;
output 	readdata_22;
output 	readdata_23;
output 	readdata_24;
output 	readdata_25;
output 	readdata_31;
output 	readdata_21;
output 	readdata_11;
output 	readdata_28;
output 	readdata_10;
output 	readdata_27;
output 	readdata_8;
output 	readdata_9;
output 	readdata_26;
output 	readdata_20;
output 	readdata_19;
output 	readdata_17;
output 	readdata_30;
output 	readdata_18;
output 	readdata_16;
output 	readdata_15;
output 	readdata_12;
output 	readdata_13;
output 	readdata_14;
output 	readdata_29;
output 	sr_0;
output 	ir_out_0;
output 	ir_out_1;
input 	d_write;
input 	r_sync_rst;
input 	W_debug_mode;
output 	oci_single_step_mode;
output 	jtag_break;
input 	saved_grant_0;
output 	waitrequest;
input 	mem_used_1;
input 	WideOr1;
input 	mem;
output 	oci_ienable_1;
output 	oci_ienable_16;
input 	[31:0] writedata_nxt;
input 	[8:0] address_nxt;
input 	debugaccess_nxt;
input 	r_early_rst;
input 	[3:0] byteenable_nxt;
input 	altera_internal_jtag;
input 	altera_internal_jtag1;
input 	state_1;
input 	state_4;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_8;
input 	splitter_nodes_receive_1_3;
input 	irf_reg_0_2;
input 	irf_reg_1_2;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[0]~q ;
wire \the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[1]~q ;
wire \the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[0] ;
wire \the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[2]~q ;
wire \the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[2]~q ;
wire \the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[1] ;
wire \the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[20]~q ;
wire \the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[20]~q ;
wire \the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[19]~q ;
wire \the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[19]~q ;
wire \the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[3]~q ;
wire \the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[2] ;
wire \the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[21]~q ;
wire \the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[21]~q ;
wire \the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[20] ;
wire \the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[19] ;
wire \the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[18]~q ;
wire \the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[17]~q ;
wire \the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[17]~q ;
wire \the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[16]~q ;
wire \the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[16]~q ;
wire \the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[24]~q ;
wire \the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[24]~q ;
wire \the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[4]~q ;
wire \the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[3] ;
wire \the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[25]~q ;
wire \the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[25]~q ;
wire \the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[26]~q ;
wire \the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[26]~q ;
wire \the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[27]~q ;
wire \the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[27]~q ;
wire \the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[22]~q ;
wire \the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[21] ;
wire \the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[18] ;
wire \the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[17] ;
wire \the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[16] ;
wire \the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[4] ;
wire \the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[5] ;
wire \the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[6] ;
wire \the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[7] ;
wire \the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[24] ;
wire \the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[5]~q ;
wire \the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[25] ;
wire \the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[26] ;
wire \the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[28]~q ;
wire \the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[28]~q ;
wire \the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[27] ;
wire \the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[29]~q ;
wire \the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[30]~q ;
wire \the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[30]~q ;
wire \the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[31]~q ;
wire \the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[31]~q ;
wire \the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[22] ;
wire \the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[23] ;
wire \the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[31] ;
wire \the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[11] ;
wire \the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[28] ;
wire \the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[10] ;
wire \the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[8] ;
wire \the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[9] ;
wire \the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[30] ;
wire \the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[15] ;
wire \the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[12] ;
wire \the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[13] ;
wire \the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[14] ;
wire \the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[29] ;
wire \the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[23]~q ;
wire \the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[23]~q ;
wire \the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[6]~q ;
wire \the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[7]~q ;
wire \the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[6]~q ;
wire \the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[11]~q ;
wire \the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[10]~q ;
wire \the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[9]~q ;
wire \the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[13]~q ;
wire \the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[14]~q ;
wire \the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[15]~q ;
wire \the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[7]~q ;
wire \the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[8]~q ;
wire \the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[9]~q ;
wire \the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[13]~q ;
wire \the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[12]~q ;
wire \the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[10]~q ;
wire \the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[11]~q ;
wire \the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[14]~q ;
wire \the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[0]~q ;
wire \writedata[3]~q ;
wire \address[0]~q ;
wire \address[3]~q ;
wire \address[2]~q ;
wire \address[1]~q ;
wire \address[7]~q ;
wire \address[6]~q ;
wire \address[5]~q ;
wire \address[4]~q ;
wire \the_first_nios2_system_cpu_cpu_nios2_avalon_reg|Equal0~1_combout ;
wire \debugaccess~q ;
wire \write~q ;
wire \the_first_nios2_system_cpu_cpu_nios2_avalon_reg|take_action_ocireg~0_combout ;
wire \the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[34]~q ;
wire \the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[35]~q ;
wire \the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|ir[1]~q ;
wire \the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|ir[0]~q ;
wire \the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|enable_action_strobe~q ;
wire \the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|take_action_ocimem_a~0_combout ;
wire \the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|take_action_ocimem_a~1_combout ;
wire \the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|take_action_ocimem_a~combout ;
wire \the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[21]~q ;
wire \the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[20]~q ;
wire \read~q ;
wire \the_first_nios2_system_cpu_cpu_nios2_oci_debug|monitor_ready~q ;
wire \the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[1]~q ;
wire \the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[0]~q ;
wire \the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[36]~q ;
wire \the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[37]~q ;
wire \the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[3]~q ;
wire \write~0_combout ;
wire \the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[19]~q ;
wire \the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[18]~q ;
wire \the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[17]~q ;
wire \read~0_combout ;
wire \the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[25]~q ;
wire \writedata[0]~q ;
wire \the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[1]~q ;
wire \the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[4]~q ;
wire \the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[26]~q ;
wire \the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[27]~q ;
wire \the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[28]~q ;
wire \byteenable[0]~q ;
wire \writedata[1]~q ;
wire \writedata[16]~q ;
wire \the_first_nios2_system_cpu_cpu_nios2_oci_debug|monitor_error~q ;
wire \the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[3]~q ;
wire \the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[2]~q ;
wire \the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[5]~q ;
wire \the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[29]~q ;
wire \the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[30]~q ;
wire \the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[31]~q ;
wire \the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[32]~q ;
wire \the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[33]~q ;
wire \the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[23]~q ;
wire \the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[22]~q ;
wire \the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[18]~q ;
wire \the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[4]~q ;
wire \the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[6]~q ;
wire \writedata[2]~q ;
wire \the_first_nios2_system_cpu_cpu_nios2_avalon_reg|oci_reg_readdata~0_combout ;
wire \the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[22]~q ;
wire \the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[24]~q ;
wire \writedata[20]~q ;
wire \byteenable[2]~q ;
wire \writedata[19]~q ;
wire \the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[16]~q ;
wire \the_first_nios2_system_cpu_cpu_nios2_avalon_reg|oci_reg_readdata[1]~1_combout ;
wire \the_first_nios2_system_cpu_cpu_nios2_oci_debug|monitor_go~q ;
wire \the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[5]~q ;
wire \the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[7]~q ;
wire \the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[29]~q ;
wire \the_first_nios2_system_cpu_cpu_nios2_oci_debug|resetlatch~q ;
wire \the_first_nios2_system_cpu_cpu_nios2_avalon_reg|oci_reg_readdata~2_combout ;
wire \writedata[21]~q ;
wire \writedata[18]~q ;
wire \writedata[17]~q ;
wire \writedata[4]~q ;
wire \writedata[5]~q ;
wire \writedata[6]~q ;
wire \writedata[7]~q ;
wire \writedata[24]~q ;
wire \byteenable[3]~q ;
wire \the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[8]~q ;
wire \writedata[25]~q ;
wire \writedata[26]~q ;
wire \writedata[27]~q ;
wire \writedata[22]~q ;
wire \writedata[23]~q ;
wire \writedata[31]~q ;
wire \writedata[11]~q ;
wire \byteenable[1]~q ;
wire \writedata[28]~q ;
wire \writedata[10]~q ;
wire \the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[8]~q ;
wire \writedata[8]~q ;
wire \writedata[9]~q ;
wire \writedata[30]~q ;
wire \the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[15]~q ;
wire \writedata[15]~q ;
wire \the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[12]~q ;
wire \writedata[12]~q ;
wire \writedata[13]~q ;
wire \writedata[14]~q ;
wire \writedata[29]~q ;
wire \the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[9]~q ;
wire \the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[10]~q ;
wire \the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[14]~q ;
wire \the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[13]~q ;
wire \the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[11]~q ;
wire \the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[12]~q ;
wire \the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[15]~q ;
wire \readdata~0_combout ;
wire \address[8]~q ;
wire \readdata~1_combout ;
wire \readdata~2_combout ;


first_nios2_system_first_nios2_system_cpu_cpu_nios2_oci_break the_first_nios2_system_cpu_cpu_nios2_oci_break(
	.break_readreg_0(\the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[0]~q ),
	.break_readreg_1(\the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[1]~q ),
	.break_readreg_2(\the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[2]~q ),
	.break_readreg_20(\the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[20]~q ),
	.break_readreg_19(\the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[19]~q ),
	.break_readreg_3(\the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[3]~q ),
	.break_readreg_21(\the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[21]~q ),
	.break_readreg_18(\the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[18]~q ),
	.break_readreg_17(\the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[17]~q ),
	.break_readreg_16(\the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[16]~q ),
	.break_readreg_24(\the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[24]~q ),
	.break_readreg_4(\the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[4]~q ),
	.break_readreg_25(\the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[25]~q ),
	.break_readreg_26(\the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[26]~q ),
	.break_readreg_27(\the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[27]~q ),
	.break_readreg_22(\the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[22]~q ),
	.break_readreg_5(\the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[5]~q ),
	.break_readreg_28(\the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[28]~q ),
	.break_readreg_29(\the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[29]~q ),
	.break_readreg_30(\the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[30]~q ),
	.break_readreg_31(\the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[31]~q ),
	.break_readreg_23(\the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[23]~q ),
	.break_readreg_6(\the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[6]~q ),
	.break_readreg_15(\the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[15]~q ),
	.break_readreg_7(\the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[7]~q ),
	.break_readreg_8(\the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[8]~q ),
	.break_readreg_9(\the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[9]~q ),
	.break_readreg_13(\the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[13]~q ),
	.break_readreg_12(\the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[12]~q ),
	.break_readreg_10(\the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[10]~q ),
	.break_readreg_11(\the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[11]~q ),
	.break_readreg_14(\the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[14]~q ),
	.ir_1(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|ir[1]~q ),
	.ir_0(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|ir[0]~q ),
	.enable_action_strobe(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|enable_action_strobe~q ),
	.jdo_21(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[21]~q ),
	.jdo_20(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[20]~q ),
	.jdo_0(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[0]~q ),
	.jdo_36(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[36]~q ),
	.jdo_37(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[37]~q ),
	.jdo_3(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[3]~q ),
	.jdo_19(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[19]~q ),
	.jdo_18(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[18]~q ),
	.jdo_17(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[17]~q ),
	.jdo_25(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[25]~q ),
	.jdo_1(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[1]~q ),
	.jdo_4(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[4]~q ),
	.jdo_26(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[26]~q ),
	.jdo_27(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[27]~q ),
	.jdo_28(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[28]~q ),
	.jdo_2(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[2]~q ),
	.jdo_5(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[5]~q ),
	.jdo_29(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[29]~q ),
	.jdo_30(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[30]~q ),
	.jdo_31(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[31]~q ),
	.jdo_23(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[23]~q ),
	.jdo_22(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[22]~q ),
	.jdo_6(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[6]~q ),
	.jdo_24(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[24]~q ),
	.jdo_16(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[16]~q ),
	.jdo_7(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[7]~q ),
	.jdo_8(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[8]~q ),
	.jdo_9(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[9]~q ),
	.jdo_10(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[10]~q ),
	.jdo_14(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[14]~q ),
	.jdo_13(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[13]~q ),
	.jdo_11(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[11]~q ),
	.jdo_12(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[12]~q ),
	.jdo_15(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[15]~q ),
	.clk_clk(clk_clk));

first_nios2_system_first_nios2_system_cpu_cpu_nios2_oci_debug the_first_nios2_system_cpu_cpu_nios2_oci_debug(
	.r_sync_rst(r_sync_rst),
	.jtag_break1(jtag_break),
	.take_action_ocireg(\the_first_nios2_system_cpu_cpu_nios2_avalon_reg|take_action_ocireg~0_combout ),
	.jdo_34(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[34]~q ),
	.jdo_35(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[35]~q ),
	.take_action_ocimem_a(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|take_action_ocimem_a~0_combout ),
	.take_action_ocimem_a1(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|take_action_ocimem_a~combout ),
	.jdo_21(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[21]~q ),
	.jdo_20(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[20]~q ),
	.monitor_ready1(\the_first_nios2_system_cpu_cpu_nios2_oci_debug|monitor_ready~q ),
	.jdo_19(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[19]~q ),
	.jdo_18(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[18]~q ),
	.jdo_25(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[25]~q ),
	.writedata_0(\writedata[0]~q ),
	.writedata_1(\writedata[1]~q ),
	.monitor_error1(\the_first_nios2_system_cpu_cpu_nios2_oci_debug|monitor_error~q ),
	.jdo_23(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[23]~q ),
	.jdo_24(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[24]~q ),
	.monitor_go1(\the_first_nios2_system_cpu_cpu_nios2_oci_debug|monitor_go~q ),
	.resetlatch1(\the_first_nios2_system_cpu_cpu_nios2_oci_debug|resetlatch~q ),
	.state_1(state_1),
	.clk_clk(clk_clk));

first_nios2_system_first_nios2_system_cpu_cpu_debug_slave_wrapper the_first_nios2_system_cpu_cpu_debug_slave_wrapper(
	.break_readreg_0(\the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[0]~q ),
	.break_readreg_1(\the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[1]~q ),
	.break_readreg_2(\the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[2]~q ),
	.MonDReg_2(\the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[2]~q ),
	.break_readreg_20(\the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[20]~q ),
	.MonDReg_20(\the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[20]~q ),
	.break_readreg_19(\the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[19]~q ),
	.MonDReg_19(\the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[19]~q ),
	.break_readreg_3(\the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[3]~q ),
	.break_readreg_21(\the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[21]~q ),
	.MonDReg_21(\the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[21]~q ),
	.break_readreg_18(\the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[18]~q ),
	.break_readreg_17(\the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[17]~q ),
	.MonDReg_17(\the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[17]~q ),
	.break_readreg_16(\the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[16]~q ),
	.MonDReg_16(\the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[16]~q ),
	.break_readreg_24(\the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[24]~q ),
	.MonDReg_24(\the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[24]~q ),
	.break_readreg_4(\the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[4]~q ),
	.break_readreg_25(\the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[25]~q ),
	.MonDReg_25(\the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[25]~q ),
	.break_readreg_26(\the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[26]~q ),
	.MonDReg_26(\the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[26]~q ),
	.break_readreg_27(\the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[27]~q ),
	.MonDReg_27(\the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[27]~q ),
	.break_readreg_22(\the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[22]~q ),
	.break_readreg_5(\the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[5]~q ),
	.break_readreg_28(\the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[28]~q ),
	.MonDReg_28(\the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[28]~q ),
	.break_readreg_29(\the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[29]~q ),
	.MonDReg_30(\the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[30]~q ),
	.break_readreg_30(\the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[30]~q ),
	.break_readreg_31(\the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[31]~q ),
	.MonDReg_31(\the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[31]~q ),
	.break_readreg_23(\the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[23]~q ),
	.MonDReg_23(\the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[23]~q ),
	.MonDReg_6(\the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[6]~q ),
	.MonDReg_7(\the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[7]~q ),
	.break_readreg_6(\the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[6]~q ),
	.MonDReg_11(\the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[11]~q ),
	.MonDReg_10(\the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[10]~q ),
	.MonDReg_9(\the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[9]~q ),
	.MonDReg_13(\the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[13]~q ),
	.MonDReg_14(\the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[14]~q ),
	.break_readreg_15(\the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[15]~q ),
	.break_readreg_7(\the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[7]~q ),
	.break_readreg_8(\the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[8]~q ),
	.break_readreg_9(\the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[9]~q ),
	.break_readreg_13(\the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[13]~q ),
	.break_readreg_12(\the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[12]~q ),
	.break_readreg_10(\the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[10]~q ),
	.break_readreg_11(\the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[11]~q ),
	.break_readreg_14(\the_first_nios2_system_cpu_cpu_nios2_oci_break|break_readreg[14]~q ),
	.sr_0(sr_0),
	.ir_out_0(ir_out_0),
	.ir_out_1(ir_out_1),
	.W_debug_mode(W_debug_mode),
	.MonDReg_0(\the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[0]~q ),
	.jdo_34(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[34]~q ),
	.jdo_35(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[35]~q ),
	.ir_1(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|ir[1]~q ),
	.ir_0(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|ir[0]~q ),
	.enable_action_strobe(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|enable_action_strobe~q ),
	.take_action_ocimem_a(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|take_action_ocimem_a~0_combout ),
	.take_action_ocimem_a1(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|take_action_ocimem_a~1_combout ),
	.take_action_ocimem_a2(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|take_action_ocimem_a~combout ),
	.jdo_21(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[21]~q ),
	.jdo_20(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[20]~q ),
	.monitor_ready(\the_first_nios2_system_cpu_cpu_nios2_oci_debug|monitor_ready~q ),
	.MonDReg_1(\the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[1]~q ),
	.jdo_0(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[0]~q ),
	.jdo_36(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[36]~q ),
	.jdo_37(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[37]~q ),
	.jdo_3(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[3]~q ),
	.jdo_19(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[19]~q ),
	.jdo_18(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[18]~q ),
	.jdo_17(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[17]~q ),
	.jdo_25(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[25]~q ),
	.jdo_1(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[1]~q ),
	.jdo_4(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[4]~q ),
	.jdo_26(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[26]~q ),
	.jdo_27(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[27]~q ),
	.jdo_28(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[28]~q ),
	.monitor_error(\the_first_nios2_system_cpu_cpu_nios2_oci_debug|monitor_error~q ),
	.MonDReg_3(\the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[3]~q ),
	.jdo_2(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[2]~q ),
	.jdo_5(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[5]~q ),
	.jdo_29(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[29]~q ),
	.jdo_30(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[30]~q ),
	.jdo_31(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[31]~q ),
	.jdo_32(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[32]~q ),
	.jdo_33(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[33]~q ),
	.jdo_23(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[23]~q ),
	.jdo_22(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[22]~q ),
	.MonDReg_18(\the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[18]~q ),
	.MonDReg_4(\the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[4]~q ),
	.jdo_6(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[6]~q ),
	.MonDReg_22(\the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[22]~q ),
	.jdo_24(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[24]~q ),
	.jdo_16(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[16]~q ),
	.MonDReg_5(\the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[5]~q ),
	.jdo_7(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[7]~q ),
	.MonDReg_29(\the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[29]~q ),
	.resetlatch(\the_first_nios2_system_cpu_cpu_nios2_oci_debug|resetlatch~q ),
	.jdo_8(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[8]~q ),
	.MonDReg_8(\the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[8]~q ),
	.MonDReg_15(\the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[15]~q ),
	.MonDReg_12(\the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[12]~q ),
	.jdo_9(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[9]~q ),
	.jdo_10(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[10]~q ),
	.jdo_14(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[14]~q ),
	.jdo_13(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[13]~q ),
	.jdo_11(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[11]~q ),
	.jdo_12(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[12]~q ),
	.jdo_15(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[15]~q ),
	.altera_internal_jtag(altera_internal_jtag),
	.altera_internal_jtag1(altera_internal_jtag1),
	.state_4(state_4),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.state_8(state_8),
	.splitter_nodes_receive_1_3(splitter_nodes_receive_1_3),
	.irf_reg_0_2(irf_reg_0_2),
	.irf_reg_1_2(irf_reg_1_2),
	.clk_clk(clk_clk));

first_nios2_system_first_nios2_system_cpu_cpu_nios2_ocimem the_first_nios2_system_cpu_cpu_nios2_ocimem(
	.q_a_0(\the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[0] ),
	.MonDReg_2(\the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[2]~q ),
	.q_a_1(\the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[1] ),
	.MonDReg_20(\the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[20]~q ),
	.MonDReg_19(\the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[19]~q ),
	.q_a_2(\the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[2] ),
	.MonDReg_21(\the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[21]~q ),
	.q_a_20(\the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[20] ),
	.q_a_19(\the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[19] ),
	.MonDReg_17(\the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[17]~q ),
	.MonDReg_16(\the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[16]~q ),
	.MonDReg_24(\the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[24]~q ),
	.q_a_3(\the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[3] ),
	.MonDReg_25(\the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[25]~q ),
	.MonDReg_26(\the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[26]~q ),
	.MonDReg_27(\the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[27]~q ),
	.q_a_21(\the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[21] ),
	.q_a_18(\the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[18] ),
	.q_a_17(\the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[17] ),
	.q_a_16(\the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[16] ),
	.q_a_4(\the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[4] ),
	.q_a_5(\the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[5] ),
	.q_a_6(\the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[6] ),
	.q_a_7(\the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[7] ),
	.q_a_24(\the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[24] ),
	.q_a_25(\the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[25] ),
	.q_a_26(\the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[26] ),
	.MonDReg_28(\the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[28]~q ),
	.q_a_27(\the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[27] ),
	.MonDReg_30(\the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[30]~q ),
	.MonDReg_31(\the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[31]~q ),
	.q_a_22(\the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[22] ),
	.q_a_23(\the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[23] ),
	.q_a_31(\the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[31] ),
	.q_a_11(\the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[11] ),
	.q_a_28(\the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[28] ),
	.q_a_10(\the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[10] ),
	.q_a_8(\the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[8] ),
	.q_a_9(\the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[9] ),
	.q_a_30(\the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[30] ),
	.q_a_15(\the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[15] ),
	.q_a_12(\the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[12] ),
	.q_a_13(\the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[13] ),
	.q_a_14(\the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[14] ),
	.q_a_29(\the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[29] ),
	.MonDReg_23(\the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[23]~q ),
	.MonDReg_6(\the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[6]~q ),
	.MonDReg_7(\the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[7]~q ),
	.MonDReg_11(\the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[11]~q ),
	.MonDReg_10(\the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[10]~q ),
	.MonDReg_9(\the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[9]~q ),
	.MonDReg_13(\the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[13]~q ),
	.MonDReg_14(\the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[14]~q ),
	.waitrequest1(waitrequest),
	.MonDReg_0(\the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[0]~q ),
	.writedata_3(\writedata[3]~q ),
	.address_0(\address[0]~q ),
	.address_3(\address[3]~q ),
	.address_2(\address[2]~q ),
	.address_1(\address[1]~q ),
	.address_8(\address[8]~q ),
	.address_7(\address[7]~q ),
	.address_6(\address[6]~q ),
	.address_5(\address[5]~q ),
	.address_4(\address[4]~q ),
	.debugaccess(\debugaccess~q ),
	.write(\write~q ),
	.jdo_34(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[34]~q ),
	.jdo_35(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[35]~q ),
	.take_action_ocimem_a(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|take_action_ocimem_a~0_combout ),
	.take_no_action_ocimem_a(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|take_action_ocimem_a~1_combout ),
	.take_action_ocimem_a1(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|take_action_ocimem_a~combout ),
	.jdo_21(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[21]~q ),
	.jdo_20(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[20]~q ),
	.read(\read~q ),
	.MonDReg_1(\the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[1]~q ),
	.jdo_3(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[3]~q ),
	.jdo_19(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[19]~q ),
	.jdo_18(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[18]~q ),
	.jdo_17(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[17]~q ),
	.jdo_25(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[25]~q ),
	.writedata_0(\writedata[0]~q ),
	.jdo_4(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[4]~q ),
	.jdo_26(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[26]~q ),
	.jdo_27(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[27]~q ),
	.jdo_28(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[28]~q ),
	.r_early_rst(r_early_rst),
	.byteenable_0(\byteenable[0]~q ),
	.writedata_1(\writedata[1]~q ),
	.writedata_16(\writedata[16]~q ),
	.MonDReg_3(\the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[3]~q ),
	.jdo_5(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[5]~q ),
	.jdo_29(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[29]~q ),
	.jdo_30(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[30]~q ),
	.jdo_31(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[31]~q ),
	.jdo_32(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[32]~q ),
	.jdo_33(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[33]~q ),
	.jdo_23(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[23]~q ),
	.jdo_22(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[22]~q ),
	.MonDReg_18(\the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[18]~q ),
	.MonDReg_4(\the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[4]~q ),
	.jdo_6(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[6]~q ),
	.writedata_2(\writedata[2]~q ),
	.MonDReg_22(\the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[22]~q ),
	.jdo_24(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[24]~q ),
	.writedata_20(\writedata[20]~q ),
	.byteenable_2(\byteenable[2]~q ),
	.writedata_19(\writedata[19]~q ),
	.jdo_16(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[16]~q ),
	.MonDReg_5(\the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[5]~q ),
	.jdo_7(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[7]~q ),
	.MonDReg_29(\the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[29]~q ),
	.writedata_21(\writedata[21]~q ),
	.writedata_18(\writedata[18]~q ),
	.writedata_17(\writedata[17]~q ),
	.writedata_4(\writedata[4]~q ),
	.writedata_5(\writedata[5]~q ),
	.writedata_6(\writedata[6]~q ),
	.writedata_7(\writedata[7]~q ),
	.writedata_24(\writedata[24]~q ),
	.byteenable_3(\byteenable[3]~q ),
	.jdo_8(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[8]~q ),
	.writedata_25(\writedata[25]~q ),
	.writedata_26(\writedata[26]~q ),
	.writedata_27(\writedata[27]~q ),
	.writedata_22(\writedata[22]~q ),
	.writedata_23(\writedata[23]~q ),
	.writedata_31(\writedata[31]~q ),
	.writedata_11(\writedata[11]~q ),
	.byteenable_1(\byteenable[1]~q ),
	.writedata_28(\writedata[28]~q ),
	.writedata_10(\writedata[10]~q ),
	.MonDReg_8(\the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[8]~q ),
	.writedata_8(\writedata[8]~q ),
	.writedata_9(\writedata[9]~q ),
	.writedata_30(\writedata[30]~q ),
	.MonDReg_15(\the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[15]~q ),
	.writedata_15(\writedata[15]~q ),
	.MonDReg_12(\the_first_nios2_system_cpu_cpu_nios2_ocimem|MonDReg[12]~q ),
	.writedata_12(\writedata[12]~q ),
	.writedata_13(\writedata[13]~q ),
	.writedata_14(\writedata[14]~q ),
	.writedata_29(\writedata[29]~q ),
	.jdo_9(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[9]~q ),
	.jdo_10(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[10]~q ),
	.jdo_14(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[14]~q ),
	.jdo_13(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[13]~q ),
	.jdo_11(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[11]~q ),
	.jdo_12(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[12]~q ),
	.jdo_15(\the_first_nios2_system_cpu_cpu_debug_slave_wrapper|the_first_nios2_system_cpu_cpu_debug_slave_sysclk|jdo[15]~q ),
	.clk_clk(clk_clk));

first_nios2_system_first_nios2_system_cpu_cpu_nios2_avalon_reg the_first_nios2_system_cpu_cpu_nios2_avalon_reg(
	.r_sync_rst(r_sync_rst),
	.oci_single_step_mode1(oci_single_step_mode),
	.writedata_3(\writedata[3]~q ),
	.address_0(\address[0]~q ),
	.address_3(\address[3]~q ),
	.address_2(\address[2]~q ),
	.address_1(\address[1]~q ),
	.address_8(\address[8]~q ),
	.address_7(\address[7]~q ),
	.address_6(\address[6]~q ),
	.address_5(\address[5]~q ),
	.address_4(\address[4]~q ),
	.Equal0(\the_first_nios2_system_cpu_cpu_nios2_avalon_reg|Equal0~1_combout ),
	.debugaccess(\debugaccess~q ),
	.write(\write~q ),
	.take_action_ocireg(\the_first_nios2_system_cpu_cpu_nios2_avalon_reg|take_action_ocireg~0_combout ),
	.monitor_ready(\the_first_nios2_system_cpu_cpu_nios2_oci_debug|monitor_ready~q ),
	.oci_ienable_1(oci_ienable_1),
	.oci_ienable_16(oci_ienable_16),
	.writedata_1(\writedata[1]~q ),
	.writedata_16(\writedata[16]~q ),
	.oci_reg_readdata(\the_first_nios2_system_cpu_cpu_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.oci_reg_readdata_1(\the_first_nios2_system_cpu_cpu_nios2_avalon_reg|oci_reg_readdata[1]~1_combout ),
	.oci_reg_readdata1(\the_first_nios2_system_cpu_cpu_nios2_avalon_reg|oci_reg_readdata~2_combout ),
	.clk_clk(clk_clk));

dffeas \writedata[3] (
	.clk(clk_clk),
	.d(writedata_nxt[3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[3]~q ),
	.prn(vcc));
defparam \writedata[3] .is_wysiwyg = "true";
defparam \writedata[3] .power_up = "low";

dffeas \address[0] (
	.clk(clk_clk),
	.d(address_nxt[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[0]~q ),
	.prn(vcc));
defparam \address[0] .is_wysiwyg = "true";
defparam \address[0] .power_up = "low";

dffeas \address[3] (
	.clk(clk_clk),
	.d(address_nxt[3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[3]~q ),
	.prn(vcc));
defparam \address[3] .is_wysiwyg = "true";
defparam \address[3] .power_up = "low";

dffeas \address[2] (
	.clk(clk_clk),
	.d(address_nxt[2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[2]~q ),
	.prn(vcc));
defparam \address[2] .is_wysiwyg = "true";
defparam \address[2] .power_up = "low";

dffeas \address[1] (
	.clk(clk_clk),
	.d(address_nxt[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[1]~q ),
	.prn(vcc));
defparam \address[1] .is_wysiwyg = "true";
defparam \address[1] .power_up = "low";

dffeas \address[7] (
	.clk(clk_clk),
	.d(address_nxt[7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[7]~q ),
	.prn(vcc));
defparam \address[7] .is_wysiwyg = "true";
defparam \address[7] .power_up = "low";

dffeas \address[6] (
	.clk(clk_clk),
	.d(address_nxt[6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[6]~q ),
	.prn(vcc));
defparam \address[6] .is_wysiwyg = "true";
defparam \address[6] .power_up = "low";

dffeas \address[5] (
	.clk(clk_clk),
	.d(address_nxt[5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[5]~q ),
	.prn(vcc));
defparam \address[5] .is_wysiwyg = "true";
defparam \address[5] .power_up = "low";

dffeas \address[4] (
	.clk(clk_clk),
	.d(address_nxt[4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[4]~q ),
	.prn(vcc));
defparam \address[4] .is_wysiwyg = "true";
defparam \address[4] .power_up = "low";

dffeas debugaccess(
	.clk(clk_clk),
	.d(debugaccess_nxt),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\debugaccess~q ),
	.prn(vcc));
defparam debugaccess.is_wysiwyg = "true";
defparam debugaccess.power_up = "low";

dffeas write(
	.clk(clk_clk),
	.d(\write~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\write~q ),
	.prn(vcc));
defparam write.is_wysiwyg = "true";
defparam write.power_up = "low";

dffeas read(
	.clk(clk_clk),
	.d(\read~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\read~q ),
	.prn(vcc));
defparam read.is_wysiwyg = "true";
defparam read.power_up = "low";

cyclonev_lcell_comb \write~0 (
	.dataa(!d_write),
	.datab(!saved_grant_0),
	.datac(!waitrequest),
	.datad(!mem_used_1),
	.datae(!\write~q ),
	.dataf(!WideOr1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\write~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \write~0 .extended_lut = "off";
defparam \write~0 .lut_mask = 64'hFF7FFFFFFF7F7F7F;
defparam \write~0 .shared_arith = "off";

cyclonev_lcell_comb \read~0 (
	.dataa(!waitrequest),
	.datab(!mem_used_1),
	.datac(!WideOr1),
	.datad(!mem),
	.datae(!\read~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read~0 .extended_lut = "off";
defparam \read~0 .lut_mask = 64'hDDFFF5FFDDFFF5FF;
defparam \read~0 .shared_arith = "off";

dffeas \writedata[0] (
	.clk(clk_clk),
	.d(writedata_nxt[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[0]~q ),
	.prn(vcc));
defparam \writedata[0] .is_wysiwyg = "true";
defparam \writedata[0] .power_up = "low";

dffeas \byteenable[0] (
	.clk(clk_clk),
	.d(byteenable_nxt[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\byteenable[0]~q ),
	.prn(vcc));
defparam \byteenable[0] .is_wysiwyg = "true";
defparam \byteenable[0] .power_up = "low";

dffeas \writedata[1] (
	.clk(clk_clk),
	.d(writedata_nxt[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[1]~q ),
	.prn(vcc));
defparam \writedata[1] .is_wysiwyg = "true";
defparam \writedata[1] .power_up = "low";

dffeas \writedata[16] (
	.clk(clk_clk),
	.d(writedata_nxt[16]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[16]~q ),
	.prn(vcc));
defparam \writedata[16] .is_wysiwyg = "true";
defparam \writedata[16] .power_up = "low";

dffeas \writedata[2] (
	.clk(clk_clk),
	.d(writedata_nxt[2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[2]~q ),
	.prn(vcc));
defparam \writedata[2] .is_wysiwyg = "true";
defparam \writedata[2] .power_up = "low";

dffeas \writedata[20] (
	.clk(clk_clk),
	.d(writedata_nxt[20]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[20]~q ),
	.prn(vcc));
defparam \writedata[20] .is_wysiwyg = "true";
defparam \writedata[20] .power_up = "low";

dffeas \byteenable[2] (
	.clk(clk_clk),
	.d(byteenable_nxt[2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\byteenable[2]~q ),
	.prn(vcc));
defparam \byteenable[2] .is_wysiwyg = "true";
defparam \byteenable[2] .power_up = "low";

dffeas \writedata[19] (
	.clk(clk_clk),
	.d(writedata_nxt[19]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[19]~q ),
	.prn(vcc));
defparam \writedata[19] .is_wysiwyg = "true";
defparam \writedata[19] .power_up = "low";

dffeas \writedata[21] (
	.clk(clk_clk),
	.d(writedata_nxt[21]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[21]~q ),
	.prn(vcc));
defparam \writedata[21] .is_wysiwyg = "true";
defparam \writedata[21] .power_up = "low";

dffeas \writedata[18] (
	.clk(clk_clk),
	.d(writedata_nxt[18]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[18]~q ),
	.prn(vcc));
defparam \writedata[18] .is_wysiwyg = "true";
defparam \writedata[18] .power_up = "low";

dffeas \writedata[17] (
	.clk(clk_clk),
	.d(writedata_nxt[17]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[17]~q ),
	.prn(vcc));
defparam \writedata[17] .is_wysiwyg = "true";
defparam \writedata[17] .power_up = "low";

dffeas \writedata[4] (
	.clk(clk_clk),
	.d(writedata_nxt[4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[4]~q ),
	.prn(vcc));
defparam \writedata[4] .is_wysiwyg = "true";
defparam \writedata[4] .power_up = "low";

dffeas \writedata[5] (
	.clk(clk_clk),
	.d(writedata_nxt[5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[5]~q ),
	.prn(vcc));
defparam \writedata[5] .is_wysiwyg = "true";
defparam \writedata[5] .power_up = "low";

dffeas \writedata[6] (
	.clk(clk_clk),
	.d(writedata_nxt[6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[6]~q ),
	.prn(vcc));
defparam \writedata[6] .is_wysiwyg = "true";
defparam \writedata[6] .power_up = "low";

dffeas \writedata[7] (
	.clk(clk_clk),
	.d(writedata_nxt[7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[7]~q ),
	.prn(vcc));
defparam \writedata[7] .is_wysiwyg = "true";
defparam \writedata[7] .power_up = "low";

dffeas \writedata[24] (
	.clk(clk_clk),
	.d(writedata_nxt[24]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[24]~q ),
	.prn(vcc));
defparam \writedata[24] .is_wysiwyg = "true";
defparam \writedata[24] .power_up = "low";

dffeas \byteenable[3] (
	.clk(clk_clk),
	.d(byteenable_nxt[3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\byteenable[3]~q ),
	.prn(vcc));
defparam \byteenable[3] .is_wysiwyg = "true";
defparam \byteenable[3] .power_up = "low";

dffeas \writedata[25] (
	.clk(clk_clk),
	.d(writedata_nxt[25]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[25]~q ),
	.prn(vcc));
defparam \writedata[25] .is_wysiwyg = "true";
defparam \writedata[25] .power_up = "low";

dffeas \writedata[26] (
	.clk(clk_clk),
	.d(writedata_nxt[26]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[26]~q ),
	.prn(vcc));
defparam \writedata[26] .is_wysiwyg = "true";
defparam \writedata[26] .power_up = "low";

dffeas \writedata[27] (
	.clk(clk_clk),
	.d(writedata_nxt[27]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[27]~q ),
	.prn(vcc));
defparam \writedata[27] .is_wysiwyg = "true";
defparam \writedata[27] .power_up = "low";

dffeas \writedata[22] (
	.clk(clk_clk),
	.d(writedata_nxt[22]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[22]~q ),
	.prn(vcc));
defparam \writedata[22] .is_wysiwyg = "true";
defparam \writedata[22] .power_up = "low";

dffeas \writedata[23] (
	.clk(clk_clk),
	.d(writedata_nxt[23]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[23]~q ),
	.prn(vcc));
defparam \writedata[23] .is_wysiwyg = "true";
defparam \writedata[23] .power_up = "low";

dffeas \writedata[31] (
	.clk(clk_clk),
	.d(writedata_nxt[31]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[31]~q ),
	.prn(vcc));
defparam \writedata[31] .is_wysiwyg = "true";
defparam \writedata[31] .power_up = "low";

dffeas \writedata[11] (
	.clk(clk_clk),
	.d(writedata_nxt[11]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[11]~q ),
	.prn(vcc));
defparam \writedata[11] .is_wysiwyg = "true";
defparam \writedata[11] .power_up = "low";

dffeas \byteenable[1] (
	.clk(clk_clk),
	.d(byteenable_nxt[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\byteenable[1]~q ),
	.prn(vcc));
defparam \byteenable[1] .is_wysiwyg = "true";
defparam \byteenable[1] .power_up = "low";

dffeas \writedata[28] (
	.clk(clk_clk),
	.d(writedata_nxt[28]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[28]~q ),
	.prn(vcc));
defparam \writedata[28] .is_wysiwyg = "true";
defparam \writedata[28] .power_up = "low";

dffeas \writedata[10] (
	.clk(clk_clk),
	.d(writedata_nxt[10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[10]~q ),
	.prn(vcc));
defparam \writedata[10] .is_wysiwyg = "true";
defparam \writedata[10] .power_up = "low";

dffeas \writedata[8] (
	.clk(clk_clk),
	.d(writedata_nxt[8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[8]~q ),
	.prn(vcc));
defparam \writedata[8] .is_wysiwyg = "true";
defparam \writedata[8] .power_up = "low";

dffeas \writedata[9] (
	.clk(clk_clk),
	.d(writedata_nxt[9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[9]~q ),
	.prn(vcc));
defparam \writedata[9] .is_wysiwyg = "true";
defparam \writedata[9] .power_up = "low";

dffeas \writedata[30] (
	.clk(clk_clk),
	.d(writedata_nxt[30]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[30]~q ),
	.prn(vcc));
defparam \writedata[30] .is_wysiwyg = "true";
defparam \writedata[30] .power_up = "low";

dffeas \writedata[15] (
	.clk(clk_clk),
	.d(writedata_nxt[15]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[15]~q ),
	.prn(vcc));
defparam \writedata[15] .is_wysiwyg = "true";
defparam \writedata[15] .power_up = "low";

dffeas \writedata[12] (
	.clk(clk_clk),
	.d(writedata_nxt[12]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[12]~q ),
	.prn(vcc));
defparam \writedata[12] .is_wysiwyg = "true";
defparam \writedata[12] .power_up = "low";

dffeas \writedata[13] (
	.clk(clk_clk),
	.d(writedata_nxt[13]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[13]~q ),
	.prn(vcc));
defparam \writedata[13] .is_wysiwyg = "true";
defparam \writedata[13] .power_up = "low";

dffeas \writedata[14] (
	.clk(clk_clk),
	.d(writedata_nxt[14]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[14]~q ),
	.prn(vcc));
defparam \writedata[14] .is_wysiwyg = "true";
defparam \writedata[14] .power_up = "low";

dffeas \writedata[29] (
	.clk(clk_clk),
	.d(writedata_nxt[29]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[29]~q ),
	.prn(vcc));
defparam \writedata[29] .is_wysiwyg = "true";
defparam \writedata[29] .power_up = "low";

dffeas \readdata[0] (
	.clk(clk_clk),
	.d(\readdata~0_combout ),
	.asdata(\the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[0] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_0),
	.prn(vcc));
defparam \readdata[0] .is_wysiwyg = "true";
defparam \readdata[0] .power_up = "low";

dffeas \readdata[1] (
	.clk(clk_clk),
	.d(\the_first_nios2_system_cpu_cpu_nios2_avalon_reg|oci_reg_readdata[1]~1_combout ),
	.asdata(\the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[1] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_1),
	.prn(vcc));
defparam \readdata[1] .is_wysiwyg = "true";
defparam \readdata[1] .power_up = "low";

dffeas \readdata[2] (
	.clk(clk_clk),
	.d(\readdata~1_combout ),
	.asdata(\the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[2] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_2),
	.prn(vcc));
defparam \readdata[2] .is_wysiwyg = "true";
defparam \readdata[2] .power_up = "low";

dffeas \readdata[3] (
	.clk(clk_clk),
	.d(\readdata~2_combout ),
	.asdata(\the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[3] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_3),
	.prn(vcc));
defparam \readdata[3] .is_wysiwyg = "true";
defparam \readdata[3] .power_up = "low";

dffeas \readdata[4] (
	.clk(clk_clk),
	.d(\the_first_nios2_system_cpu_cpu_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[4] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_4),
	.prn(vcc));
defparam \readdata[4] .is_wysiwyg = "true";
defparam \readdata[4] .power_up = "low";

dffeas \readdata[5] (
	.clk(clk_clk),
	.d(\the_first_nios2_system_cpu_cpu_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[5] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_5),
	.prn(vcc));
defparam \readdata[5] .is_wysiwyg = "true";
defparam \readdata[5] .power_up = "low";

dffeas \readdata[6] (
	.clk(clk_clk),
	.d(\the_first_nios2_system_cpu_cpu_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[6] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_6),
	.prn(vcc));
defparam \readdata[6] .is_wysiwyg = "true";
defparam \readdata[6] .power_up = "low";

dffeas \readdata[7] (
	.clk(clk_clk),
	.d(\the_first_nios2_system_cpu_cpu_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[7] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_7),
	.prn(vcc));
defparam \readdata[7] .is_wysiwyg = "true";
defparam \readdata[7] .power_up = "low";

dffeas \readdata[22] (
	.clk(clk_clk),
	.d(\the_first_nios2_system_cpu_cpu_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[22] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_22),
	.prn(vcc));
defparam \readdata[22] .is_wysiwyg = "true";
defparam \readdata[22] .power_up = "low";

dffeas \readdata[23] (
	.clk(clk_clk),
	.d(\the_first_nios2_system_cpu_cpu_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[23] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_23),
	.prn(vcc));
defparam \readdata[23] .is_wysiwyg = "true";
defparam \readdata[23] .power_up = "low";

dffeas \readdata[24] (
	.clk(clk_clk),
	.d(\the_first_nios2_system_cpu_cpu_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[24] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_24),
	.prn(vcc));
defparam \readdata[24] .is_wysiwyg = "true";
defparam \readdata[24] .power_up = "low";

dffeas \readdata[25] (
	.clk(clk_clk),
	.d(\the_first_nios2_system_cpu_cpu_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[25] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_25),
	.prn(vcc));
defparam \readdata[25] .is_wysiwyg = "true";
defparam \readdata[25] .power_up = "low";

dffeas \readdata[31] (
	.clk(clk_clk),
	.d(\the_first_nios2_system_cpu_cpu_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[31] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_31),
	.prn(vcc));
defparam \readdata[31] .is_wysiwyg = "true";
defparam \readdata[31] .power_up = "low";

dffeas \readdata[21] (
	.clk(clk_clk),
	.d(\the_first_nios2_system_cpu_cpu_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[21] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_21),
	.prn(vcc));
defparam \readdata[21] .is_wysiwyg = "true";
defparam \readdata[21] .power_up = "low";

dffeas \readdata[11] (
	.clk(clk_clk),
	.d(\the_first_nios2_system_cpu_cpu_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[11] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_11),
	.prn(vcc));
defparam \readdata[11] .is_wysiwyg = "true";
defparam \readdata[11] .power_up = "low";

dffeas \readdata[28] (
	.clk(clk_clk),
	.d(\the_first_nios2_system_cpu_cpu_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[28] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_28),
	.prn(vcc));
defparam \readdata[28] .is_wysiwyg = "true";
defparam \readdata[28] .power_up = "low";

dffeas \readdata[10] (
	.clk(clk_clk),
	.d(\the_first_nios2_system_cpu_cpu_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[10] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_10),
	.prn(vcc));
defparam \readdata[10] .is_wysiwyg = "true";
defparam \readdata[10] .power_up = "low";

dffeas \readdata[27] (
	.clk(clk_clk),
	.d(\the_first_nios2_system_cpu_cpu_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[27] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_27),
	.prn(vcc));
defparam \readdata[27] .is_wysiwyg = "true";
defparam \readdata[27] .power_up = "low";

dffeas \readdata[8] (
	.clk(clk_clk),
	.d(\the_first_nios2_system_cpu_cpu_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[8] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_8),
	.prn(vcc));
defparam \readdata[8] .is_wysiwyg = "true";
defparam \readdata[8] .power_up = "low";

dffeas \readdata[9] (
	.clk(clk_clk),
	.d(\the_first_nios2_system_cpu_cpu_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[9] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_9),
	.prn(vcc));
defparam \readdata[9] .is_wysiwyg = "true";
defparam \readdata[9] .power_up = "low";

dffeas \readdata[26] (
	.clk(clk_clk),
	.d(\the_first_nios2_system_cpu_cpu_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[26] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_26),
	.prn(vcc));
defparam \readdata[26] .is_wysiwyg = "true";
defparam \readdata[26] .power_up = "low";

dffeas \readdata[20] (
	.clk(clk_clk),
	.d(\the_first_nios2_system_cpu_cpu_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[20] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_20),
	.prn(vcc));
defparam \readdata[20] .is_wysiwyg = "true";
defparam \readdata[20] .power_up = "low";

dffeas \readdata[19] (
	.clk(clk_clk),
	.d(\the_first_nios2_system_cpu_cpu_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[19] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_19),
	.prn(vcc));
defparam \readdata[19] .is_wysiwyg = "true";
defparam \readdata[19] .power_up = "low";

dffeas \readdata[17] (
	.clk(clk_clk),
	.d(\the_first_nios2_system_cpu_cpu_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[17] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_17),
	.prn(vcc));
defparam \readdata[17] .is_wysiwyg = "true";
defparam \readdata[17] .power_up = "low";

dffeas \readdata[30] (
	.clk(clk_clk),
	.d(\the_first_nios2_system_cpu_cpu_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[30] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_30),
	.prn(vcc));
defparam \readdata[30] .is_wysiwyg = "true";
defparam \readdata[30] .power_up = "low";

dffeas \readdata[18] (
	.clk(clk_clk),
	.d(\the_first_nios2_system_cpu_cpu_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[18] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_18),
	.prn(vcc));
defparam \readdata[18] .is_wysiwyg = "true";
defparam \readdata[18] .power_up = "low";

dffeas \readdata[16] (
	.clk(clk_clk),
	.d(\the_first_nios2_system_cpu_cpu_nios2_avalon_reg|oci_reg_readdata~2_combout ),
	.asdata(\the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[16] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_16),
	.prn(vcc));
defparam \readdata[16] .is_wysiwyg = "true";
defparam \readdata[16] .power_up = "low";

dffeas \readdata[15] (
	.clk(clk_clk),
	.d(\the_first_nios2_system_cpu_cpu_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[15] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_15),
	.prn(vcc));
defparam \readdata[15] .is_wysiwyg = "true";
defparam \readdata[15] .power_up = "low";

dffeas \readdata[12] (
	.clk(clk_clk),
	.d(\the_first_nios2_system_cpu_cpu_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[12] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_12),
	.prn(vcc));
defparam \readdata[12] .is_wysiwyg = "true";
defparam \readdata[12] .power_up = "low";

dffeas \readdata[13] (
	.clk(clk_clk),
	.d(\the_first_nios2_system_cpu_cpu_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[13] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_13),
	.prn(vcc));
defparam \readdata[13] .is_wysiwyg = "true";
defparam \readdata[13] .power_up = "low";

dffeas \readdata[14] (
	.clk(clk_clk),
	.d(\the_first_nios2_system_cpu_cpu_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[14] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_14),
	.prn(vcc));
defparam \readdata[14] .is_wysiwyg = "true";
defparam \readdata[14] .power_up = "low";

dffeas \readdata[29] (
	.clk(clk_clk),
	.d(\the_first_nios2_system_cpu_cpu_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[29] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_29),
	.prn(vcc));
defparam \readdata[29] .is_wysiwyg = "true";
defparam \readdata[29] .power_up = "low";

cyclonev_lcell_comb \readdata~0 (
	.dataa(!\the_first_nios2_system_cpu_cpu_nios2_avalon_reg|Equal0~1_combout ),
	.datab(!\the_first_nios2_system_cpu_cpu_nios2_oci_debug|monitor_error~q ),
	.datac(!\the_first_nios2_system_cpu_cpu_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\readdata~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata~0 .extended_lut = "off";
defparam \readdata~0 .lut_mask = 64'h2727272727272727;
defparam \readdata~0 .shared_arith = "off";

dffeas \address[8] (
	.clk(clk_clk),
	.d(address_nxt[8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[8]~q ),
	.prn(vcc));
defparam \address[8] .is_wysiwyg = "true";
defparam \address[8] .power_up = "low";

cyclonev_lcell_comb \readdata~1 (
	.dataa(!\the_first_nios2_system_cpu_cpu_nios2_avalon_reg|Equal0~1_combout ),
	.datab(!\the_first_nios2_system_cpu_cpu_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.datac(!\the_first_nios2_system_cpu_cpu_nios2_oci_debug|monitor_go~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\readdata~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata~1 .extended_lut = "off";
defparam \readdata~1 .lut_mask = 64'h2727272727272727;
defparam \readdata~1 .shared_arith = "off";

cyclonev_lcell_comb \readdata~2 (
	.dataa(!oci_single_step_mode),
	.datab(!\the_first_nios2_system_cpu_cpu_nios2_avalon_reg|Equal0~1_combout ),
	.datac(!\the_first_nios2_system_cpu_cpu_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\readdata~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata~2 .extended_lut = "off";
defparam \readdata~2 .lut_mask = 64'h4747474747474747;
defparam \readdata~2 .shared_arith = "off";

endmodule

module first_nios2_system_first_nios2_system_cpu_cpu_debug_slave_wrapper (
	break_readreg_0,
	break_readreg_1,
	break_readreg_2,
	MonDReg_2,
	break_readreg_20,
	MonDReg_20,
	break_readreg_19,
	MonDReg_19,
	break_readreg_3,
	break_readreg_21,
	MonDReg_21,
	break_readreg_18,
	break_readreg_17,
	MonDReg_17,
	break_readreg_16,
	MonDReg_16,
	break_readreg_24,
	MonDReg_24,
	break_readreg_4,
	break_readreg_25,
	MonDReg_25,
	break_readreg_26,
	MonDReg_26,
	break_readreg_27,
	MonDReg_27,
	break_readreg_22,
	break_readreg_5,
	break_readreg_28,
	MonDReg_28,
	break_readreg_29,
	MonDReg_30,
	break_readreg_30,
	break_readreg_31,
	MonDReg_31,
	break_readreg_23,
	MonDReg_23,
	MonDReg_6,
	MonDReg_7,
	break_readreg_6,
	MonDReg_11,
	MonDReg_10,
	MonDReg_9,
	MonDReg_13,
	MonDReg_14,
	break_readreg_15,
	break_readreg_7,
	break_readreg_8,
	break_readreg_9,
	break_readreg_13,
	break_readreg_12,
	break_readreg_10,
	break_readreg_11,
	break_readreg_14,
	sr_0,
	ir_out_0,
	ir_out_1,
	W_debug_mode,
	MonDReg_0,
	jdo_34,
	jdo_35,
	ir_1,
	ir_0,
	enable_action_strobe,
	take_action_ocimem_a,
	take_action_ocimem_a1,
	take_action_ocimem_a2,
	jdo_21,
	jdo_20,
	monitor_ready,
	MonDReg_1,
	jdo_0,
	jdo_36,
	jdo_37,
	jdo_3,
	jdo_19,
	jdo_18,
	jdo_17,
	jdo_25,
	jdo_1,
	jdo_4,
	jdo_26,
	jdo_27,
	jdo_28,
	monitor_error,
	MonDReg_3,
	jdo_2,
	jdo_5,
	jdo_29,
	jdo_30,
	jdo_31,
	jdo_32,
	jdo_33,
	jdo_23,
	jdo_22,
	MonDReg_18,
	MonDReg_4,
	jdo_6,
	MonDReg_22,
	jdo_24,
	jdo_16,
	MonDReg_5,
	jdo_7,
	MonDReg_29,
	resetlatch,
	jdo_8,
	MonDReg_8,
	MonDReg_15,
	MonDReg_12,
	jdo_9,
	jdo_10,
	jdo_14,
	jdo_13,
	jdo_11,
	jdo_12,
	jdo_15,
	altera_internal_jtag,
	altera_internal_jtag1,
	state_4,
	virtual_ir_scan_reg,
	state_3,
	state_8,
	splitter_nodes_receive_1_3,
	irf_reg_0_2,
	irf_reg_1_2,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	break_readreg_0;
input 	break_readreg_1;
input 	break_readreg_2;
input 	MonDReg_2;
input 	break_readreg_20;
input 	MonDReg_20;
input 	break_readreg_19;
input 	MonDReg_19;
input 	break_readreg_3;
input 	break_readreg_21;
input 	MonDReg_21;
input 	break_readreg_18;
input 	break_readreg_17;
input 	MonDReg_17;
input 	break_readreg_16;
input 	MonDReg_16;
input 	break_readreg_24;
input 	MonDReg_24;
input 	break_readreg_4;
input 	break_readreg_25;
input 	MonDReg_25;
input 	break_readreg_26;
input 	MonDReg_26;
input 	break_readreg_27;
input 	MonDReg_27;
input 	break_readreg_22;
input 	break_readreg_5;
input 	break_readreg_28;
input 	MonDReg_28;
input 	break_readreg_29;
input 	MonDReg_30;
input 	break_readreg_30;
input 	break_readreg_31;
input 	MonDReg_31;
input 	break_readreg_23;
input 	MonDReg_23;
input 	MonDReg_6;
input 	MonDReg_7;
input 	break_readreg_6;
input 	MonDReg_11;
input 	MonDReg_10;
input 	MonDReg_9;
input 	MonDReg_13;
input 	MonDReg_14;
input 	break_readreg_15;
input 	break_readreg_7;
input 	break_readreg_8;
input 	break_readreg_9;
input 	break_readreg_13;
input 	break_readreg_12;
input 	break_readreg_10;
input 	break_readreg_11;
input 	break_readreg_14;
output 	sr_0;
output 	ir_out_0;
output 	ir_out_1;
input 	W_debug_mode;
input 	MonDReg_0;
output 	jdo_34;
output 	jdo_35;
output 	ir_1;
output 	ir_0;
output 	enable_action_strobe;
output 	take_action_ocimem_a;
output 	take_action_ocimem_a1;
output 	take_action_ocimem_a2;
output 	jdo_21;
output 	jdo_20;
input 	monitor_ready;
input 	MonDReg_1;
output 	jdo_0;
output 	jdo_36;
output 	jdo_37;
output 	jdo_3;
output 	jdo_19;
output 	jdo_18;
output 	jdo_17;
output 	jdo_25;
output 	jdo_1;
output 	jdo_4;
output 	jdo_26;
output 	jdo_27;
output 	jdo_28;
input 	monitor_error;
input 	MonDReg_3;
output 	jdo_2;
output 	jdo_5;
output 	jdo_29;
output 	jdo_30;
output 	jdo_31;
output 	jdo_32;
output 	jdo_33;
output 	jdo_23;
output 	jdo_22;
input 	MonDReg_18;
input 	MonDReg_4;
output 	jdo_6;
input 	MonDReg_22;
output 	jdo_24;
output 	jdo_16;
input 	MonDReg_5;
output 	jdo_7;
input 	MonDReg_29;
input 	resetlatch;
output 	jdo_8;
input 	MonDReg_8;
input 	MonDReg_15;
input 	MonDReg_12;
output 	jdo_9;
output 	jdo_10;
output 	jdo_14;
output 	jdo_13;
output 	jdo_11;
output 	jdo_12;
output 	jdo_15;
input 	altera_internal_jtag;
input 	altera_internal_jtag1;
input 	state_4;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_8;
input 	splitter_nodes_receive_1_3;
input 	irf_reg_0_2;
input 	irf_reg_1_2;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[1]~q ;
wire \the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[2]~q ;
wire \the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[3]~q ;
wire \the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[21]~q ;
wire \the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[20]~q ;
wire \the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[4]~q ;
wire \the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[22]~q ;
wire \the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[19]~q ;
wire \the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[18]~q ;
wire \the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[17]~q ;
wire \the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[25]~q ;
wire \the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[5]~q ;
wire \the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[26]~q ;
wire \the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[27]~q ;
wire \the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[28]~q ;
wire \the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[23]~q ;
wire \the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[6]~q ;
wire \the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[29]~q ;
wire \the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[30]~q ;
wire \the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[32]~q ;
wire \the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[24]~q ;
wire \the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[16]~q ;
wire \the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[8]~q ;
wire \the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[9]~q ;
wire \the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[10]~q ;
wire \the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[14]~q ;
wire \the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[13]~q ;
wire \the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[11]~q ;
wire \the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[12]~q ;
wire \first_nios2_system_cpu_cpu_debug_slave_phy|virtual_state_sdr~0_combout ;
wire \first_nios2_system_cpu_cpu_debug_slave_phy|virtual_state_uir~combout ;
wire \the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[34]~q ;
wire \the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[35]~q ;
wire \the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[36]~q ;
wire \the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[37]~q ;
wire \first_nios2_system_cpu_cpu_debug_slave_phy|virtual_state_cdr~combout ;
wire \the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[31]~q ;
wire \the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[33]~q ;
wire \first_nios2_system_cpu_cpu_debug_slave_phy|virtual_state_udr~0_combout ;
wire \the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[7]~q ;
wire \the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[15]~q ;


first_nios2_system_sld_virtual_jtag_basic_1 first_nios2_system_cpu_cpu_debug_slave_phy(
	.virtual_state_sdr(\first_nios2_system_cpu_cpu_debug_slave_phy|virtual_state_sdr~0_combout ),
	.virtual_state_uir1(\first_nios2_system_cpu_cpu_debug_slave_phy|virtual_state_uir~combout ),
	.virtual_state_cdr1(\first_nios2_system_cpu_cpu_debug_slave_phy|virtual_state_cdr~combout ),
	.virtual_state_udr(\first_nios2_system_cpu_cpu_debug_slave_phy|virtual_state_udr~0_combout ),
	.state_4(state_4),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.state_8(state_8),
	.splitter_nodes_receive_1_3(splitter_nodes_receive_1_3));

first_nios2_system_first_nios2_system_cpu_cpu_debug_slave_sysclk the_first_nios2_system_cpu_cpu_debug_slave_sysclk(
	.sr_1(\the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[1]~q ),
	.sr_2(\the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[2]~q ),
	.sr_3(\the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[3]~q ),
	.sr_21(\the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[21]~q ),
	.sr_20(\the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[20]~q ),
	.sr_4(\the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[4]~q ),
	.sr_22(\the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[22]~q ),
	.sr_19(\the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[19]~q ),
	.sr_18(\the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[18]~q ),
	.sr_17(\the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[17]~q ),
	.sr_25(\the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[25]~q ),
	.sr_5(\the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[5]~q ),
	.sr_26(\the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[26]~q ),
	.sr_27(\the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[27]~q ),
	.sr_28(\the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[28]~q ),
	.sr_23(\the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[23]~q ),
	.sr_6(\the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[6]~q ),
	.sr_29(\the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[29]~q ),
	.sr_30(\the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[30]~q ),
	.sr_32(\the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[32]~q ),
	.sr_24(\the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[24]~q ),
	.sr_16(\the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[16]~q ),
	.sr_8(\the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[8]~q ),
	.sr_9(\the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[9]~q ),
	.sr_10(\the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[10]~q ),
	.sr_14(\the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[14]~q ),
	.sr_13(\the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[13]~q ),
	.sr_11(\the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[11]~q ),
	.sr_12(\the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[12]~q ),
	.sr_0(sr_0),
	.virtual_state_uir(\first_nios2_system_cpu_cpu_debug_slave_phy|virtual_state_uir~combout ),
	.jdo_34(jdo_34),
	.jdo_35(jdo_35),
	.ir_1(ir_1),
	.ir_0(ir_0),
	.enable_action_strobe1(enable_action_strobe),
	.take_action_ocimem_a1(take_action_ocimem_a),
	.take_action_ocimem_a2(take_action_ocimem_a1),
	.take_action_ocimem_a3(take_action_ocimem_a2),
	.jdo_21(jdo_21),
	.jdo_20(jdo_20),
	.jdo_0(jdo_0),
	.jdo_36(jdo_36),
	.jdo_37(jdo_37),
	.jdo_3(jdo_3),
	.sr_34(\the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[34]~q ),
	.sr_35(\the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[35]~q ),
	.jdo_19(jdo_19),
	.jdo_18(jdo_18),
	.jdo_17(jdo_17),
	.jdo_25(jdo_25),
	.jdo_1(jdo_1),
	.jdo_4(jdo_4),
	.sr_36(\the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[36]~q ),
	.sr_37(\the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[37]~q ),
	.jdo_26(jdo_26),
	.jdo_27(jdo_27),
	.jdo_28(jdo_28),
	.jdo_2(jdo_2),
	.jdo_5(jdo_5),
	.jdo_29(jdo_29),
	.jdo_30(jdo_30),
	.jdo_31(jdo_31),
	.jdo_32(jdo_32),
	.jdo_33(jdo_33),
	.jdo_23(jdo_23),
	.jdo_22(jdo_22),
	.jdo_6(jdo_6),
	.sr_31(\the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[31]~q ),
	.sr_33(\the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[33]~q ),
	.virtual_state_udr(\first_nios2_system_cpu_cpu_debug_slave_phy|virtual_state_udr~0_combout ),
	.jdo_24(jdo_24),
	.jdo_16(jdo_16),
	.sr_7(\the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[7]~q ),
	.jdo_7(jdo_7),
	.jdo_8(jdo_8),
	.jdo_9(jdo_9),
	.jdo_10(jdo_10),
	.jdo_14(jdo_14),
	.jdo_13(jdo_13),
	.jdo_11(jdo_11),
	.jdo_12(jdo_12),
	.jdo_15(jdo_15),
	.sr_15(\the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[15]~q ),
	.ir_in({irf_reg_1_2,irf_reg_0_2}),
	.clk_clk(clk_clk));

first_nios2_system_first_nios2_system_cpu_cpu_debug_slave_tck the_first_nios2_system_cpu_cpu_debug_slave_tck(
	.sr_1(\the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[1]~q ),
	.sr_2(\the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[2]~q ),
	.break_readreg_0(break_readreg_0),
	.sr_3(\the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[3]~q ),
	.break_readreg_1(break_readreg_1),
	.sr_21(\the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[21]~q ),
	.sr_20(\the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[20]~q ),
	.sr_4(\the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[4]~q ),
	.break_readreg_2(break_readreg_2),
	.MonDReg_2(MonDReg_2),
	.sr_22(\the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[22]~q ),
	.break_readreg_20(break_readreg_20),
	.MonDReg_20(MonDReg_20),
	.break_readreg_19(break_readreg_19),
	.MonDReg_19(MonDReg_19),
	.sr_19(\the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[19]~q ),
	.sr_18(\the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[18]~q ),
	.sr_17(\the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[17]~q ),
	.sr_25(\the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[25]~q ),
	.sr_5(\the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[5]~q ),
	.break_readreg_3(break_readreg_3),
	.sr_26(\the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[26]~q ),
	.sr_27(\the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[27]~q ),
	.sr_28(\the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[28]~q ),
	.sr_23(\the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[23]~q ),
	.break_readreg_21(break_readreg_21),
	.MonDReg_21(MonDReg_21),
	.break_readreg_18(break_readreg_18),
	.break_readreg_17(break_readreg_17),
	.MonDReg_17(MonDReg_17),
	.break_readreg_16(break_readreg_16),
	.MonDReg_16(MonDReg_16),
	.break_readreg_24(break_readreg_24),
	.MonDReg_24(MonDReg_24),
	.sr_6(\the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[6]~q ),
	.break_readreg_4(break_readreg_4),
	.break_readreg_25(break_readreg_25),
	.MonDReg_25(MonDReg_25),
	.break_readreg_26(break_readreg_26),
	.MonDReg_26(MonDReg_26),
	.sr_29(\the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[29]~q ),
	.break_readreg_27(break_readreg_27),
	.MonDReg_27(MonDReg_27),
	.sr_30(\the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[30]~q ),
	.sr_32(\the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[32]~q ),
	.sr_24(\the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[24]~q ),
	.break_readreg_22(break_readreg_22),
	.break_readreg_5(break_readreg_5),
	.break_readreg_28(break_readreg_28),
	.MonDReg_28(MonDReg_28),
	.break_readreg_29(break_readreg_29),
	.MonDReg_30(MonDReg_30),
	.break_readreg_30(break_readreg_30),
	.break_readreg_31(break_readreg_31),
	.MonDReg_31(MonDReg_31),
	.break_readreg_23(break_readreg_23),
	.MonDReg_23(MonDReg_23),
	.sr_16(\the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[16]~q ),
	.MonDReg_6(MonDReg_6),
	.MonDReg_7(MonDReg_7),
	.sr_8(\the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[8]~q ),
	.break_readreg_6(break_readreg_6),
	.MonDReg_11(MonDReg_11),
	.MonDReg_10(MonDReg_10),
	.MonDReg_9(MonDReg_9),
	.MonDReg_13(MonDReg_13),
	.MonDReg_14(MonDReg_14),
	.break_readreg_15(break_readreg_15),
	.sr_9(\the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[9]~q ),
	.break_readreg_7(break_readreg_7),
	.sr_10(\the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[10]~q ),
	.break_readreg_8(break_readreg_8),
	.sr_14(\the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[14]~q ),
	.sr_13(\the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[13]~q ),
	.sr_11(\the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[11]~q ),
	.sr_12(\the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[12]~q ),
	.break_readreg_9(break_readreg_9),
	.break_readreg_13(break_readreg_13),
	.break_readreg_12(break_readreg_12),
	.break_readreg_10(break_readreg_10),
	.break_readreg_11(break_readreg_11),
	.break_readreg_14(break_readreg_14),
	.sr_0(sr_0),
	.ir_out_0(ir_out_0),
	.ir_out_1(ir_out_1),
	.virtual_state_sdr(\first_nios2_system_cpu_cpu_debug_slave_phy|virtual_state_sdr~0_combout ),
	.W_debug_mode(W_debug_mode),
	.MonDReg_0(MonDReg_0),
	.virtual_state_uir(\first_nios2_system_cpu_cpu_debug_slave_phy|virtual_state_uir~combout ),
	.monitor_ready(monitor_ready),
	.MonDReg_1(MonDReg_1),
	.sr_34(\the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[34]~q ),
	.sr_35(\the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[35]~q ),
	.sr_36(\the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[36]~q ),
	.sr_37(\the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[37]~q ),
	.monitor_error(monitor_error),
	.virtual_state_cdr(\first_nios2_system_cpu_cpu_debug_slave_phy|virtual_state_cdr~combout ),
	.MonDReg_3(MonDReg_3),
	.MonDReg_18(MonDReg_18),
	.MonDReg_4(MonDReg_4),
	.sr_31(\the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[31]~q ),
	.sr_33(\the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[33]~q ),
	.MonDReg_22(MonDReg_22),
	.sr_7(\the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[7]~q ),
	.MonDReg_5(MonDReg_5),
	.MonDReg_29(MonDReg_29),
	.resetlatch(resetlatch),
	.MonDReg_8(MonDReg_8),
	.MonDReg_15(MonDReg_15),
	.MonDReg_12(MonDReg_12),
	.sr_15(\the_first_nios2_system_cpu_cpu_debug_slave_tck|sr[15]~q ),
	.altera_internal_jtag(altera_internal_jtag),
	.altera_internal_jtag1(altera_internal_jtag1),
	.state_4(state_4),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.splitter_nodes_receive_1_3(splitter_nodes_receive_1_3),
	.irf_reg_0_2(irf_reg_0_2),
	.irf_reg_1_2(irf_reg_1_2));

endmodule

module first_nios2_system_first_nios2_system_cpu_cpu_debug_slave_sysclk (
	sr_1,
	sr_2,
	sr_3,
	sr_21,
	sr_20,
	sr_4,
	sr_22,
	sr_19,
	sr_18,
	sr_17,
	sr_25,
	sr_5,
	sr_26,
	sr_27,
	sr_28,
	sr_23,
	sr_6,
	sr_29,
	sr_30,
	sr_32,
	sr_24,
	sr_16,
	sr_8,
	sr_9,
	sr_10,
	sr_14,
	sr_13,
	sr_11,
	sr_12,
	sr_0,
	virtual_state_uir,
	jdo_34,
	jdo_35,
	ir_1,
	ir_0,
	enable_action_strobe1,
	take_action_ocimem_a1,
	take_action_ocimem_a2,
	take_action_ocimem_a3,
	jdo_21,
	jdo_20,
	jdo_0,
	jdo_36,
	jdo_37,
	jdo_3,
	sr_34,
	sr_35,
	jdo_19,
	jdo_18,
	jdo_17,
	jdo_25,
	jdo_1,
	jdo_4,
	sr_36,
	sr_37,
	jdo_26,
	jdo_27,
	jdo_28,
	jdo_2,
	jdo_5,
	jdo_29,
	jdo_30,
	jdo_31,
	jdo_32,
	jdo_33,
	jdo_23,
	jdo_22,
	jdo_6,
	sr_31,
	sr_33,
	virtual_state_udr,
	jdo_24,
	jdo_16,
	sr_7,
	jdo_7,
	jdo_8,
	jdo_9,
	jdo_10,
	jdo_14,
	jdo_13,
	jdo_11,
	jdo_12,
	jdo_15,
	sr_15,
	ir_in,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	sr_1;
input 	sr_2;
input 	sr_3;
input 	sr_21;
input 	sr_20;
input 	sr_4;
input 	sr_22;
input 	sr_19;
input 	sr_18;
input 	sr_17;
input 	sr_25;
input 	sr_5;
input 	sr_26;
input 	sr_27;
input 	sr_28;
input 	sr_23;
input 	sr_6;
input 	sr_29;
input 	sr_30;
input 	sr_32;
input 	sr_24;
input 	sr_16;
input 	sr_8;
input 	sr_9;
input 	sr_10;
input 	sr_14;
input 	sr_13;
input 	sr_11;
input 	sr_12;
input 	sr_0;
input 	virtual_state_uir;
output 	jdo_34;
output 	jdo_35;
output 	ir_1;
output 	ir_0;
output 	enable_action_strobe1;
output 	take_action_ocimem_a1;
output 	take_action_ocimem_a2;
output 	take_action_ocimem_a3;
output 	jdo_21;
output 	jdo_20;
output 	jdo_0;
output 	jdo_36;
output 	jdo_37;
output 	jdo_3;
input 	sr_34;
input 	sr_35;
output 	jdo_19;
output 	jdo_18;
output 	jdo_17;
output 	jdo_25;
output 	jdo_1;
output 	jdo_4;
input 	sr_36;
input 	sr_37;
output 	jdo_26;
output 	jdo_27;
output 	jdo_28;
output 	jdo_2;
output 	jdo_5;
output 	jdo_29;
output 	jdo_30;
output 	jdo_31;
output 	jdo_32;
output 	jdo_33;
output 	jdo_23;
output 	jdo_22;
output 	jdo_6;
input 	sr_31;
input 	sr_33;
input 	virtual_state_udr;
output 	jdo_24;
output 	jdo_16;
input 	sr_7;
output 	jdo_7;
output 	jdo_8;
output 	jdo_9;
output 	jdo_10;
output 	jdo_14;
output 	jdo_13;
output 	jdo_11;
output 	jdo_12;
output 	jdo_15;
input 	sr_15;
input 	[1:0] ir_in;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \the_altera_std_synchronizer3|dreg[0]~q ;
wire \the_altera_std_synchronizer4|dreg[0]~q ;
wire \sync2_udr~q ;
wire \update_jdo_strobe~0_combout ;
wire \update_jdo_strobe~q ;
wire \sync2_uir~q ;
wire \jxuir~0_combout ;
wire \jxuir~q ;


first_nios2_system_altera_std_synchronizer_1 the_altera_std_synchronizer4(
	.din(virtual_state_uir),
	.dreg_0(\the_altera_std_synchronizer4|dreg[0]~q ),
	.clk(clk_clk));

first_nios2_system_altera_std_synchronizer the_altera_std_synchronizer3(
	.dreg_0(\the_altera_std_synchronizer3|dreg[0]~q ),
	.din(virtual_state_udr),
	.clk(clk_clk));

dffeas \jdo[34] (
	.clk(clk_clk),
	.d(sr_34),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_34),
	.prn(vcc));
defparam \jdo[34] .is_wysiwyg = "true";
defparam \jdo[34] .power_up = "low";

dffeas \jdo[35] (
	.clk(clk_clk),
	.d(sr_35),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_35),
	.prn(vcc));
defparam \jdo[35] .is_wysiwyg = "true";
defparam \jdo[35] .power_up = "low";

dffeas \ir[1] (
	.clk(clk_clk),
	.d(ir_in[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\jxuir~q ),
	.q(ir_1),
	.prn(vcc));
defparam \ir[1] .is_wysiwyg = "true";
defparam \ir[1] .power_up = "low";

dffeas \ir[0] (
	.clk(clk_clk),
	.d(ir_in[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\jxuir~q ),
	.q(ir_0),
	.prn(vcc));
defparam \ir[0] .is_wysiwyg = "true";
defparam \ir[0] .power_up = "low";

dffeas enable_action_strobe(
	.clk(clk_clk),
	.d(\update_jdo_strobe~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(enable_action_strobe1),
	.prn(vcc));
defparam enable_action_strobe.is_wysiwyg = "true";
defparam enable_action_strobe.power_up = "low";

cyclonev_lcell_comb \take_action_ocimem_a~0 (
	.dataa(!ir_1),
	.datab(!ir_0),
	.datac(!enable_action_strobe1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(take_action_ocimem_a1),
	.sumout(),
	.cout(),
	.shareout());
defparam \take_action_ocimem_a~0 .extended_lut = "off";
defparam \take_action_ocimem_a~0 .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \take_action_ocimem_a~0 .shared_arith = "off";

cyclonev_lcell_comb \take_action_ocimem_a~1 (
	.dataa(!jdo_35),
	.datab(!take_action_ocimem_a1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(take_action_ocimem_a2),
	.sumout(),
	.cout(),
	.shareout());
defparam \take_action_ocimem_a~1 .extended_lut = "off";
defparam \take_action_ocimem_a~1 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \take_action_ocimem_a~1 .shared_arith = "off";

cyclonev_lcell_comb take_action_ocimem_a(
	.dataa(!jdo_34),
	.datab(!take_action_ocimem_a2),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(take_action_ocimem_a3),
	.sumout(),
	.cout(),
	.shareout());
defparam take_action_ocimem_a.extended_lut = "off";
defparam take_action_ocimem_a.lut_mask = 64'h7777777777777777;
defparam take_action_ocimem_a.shared_arith = "off";

dffeas \jdo[21] (
	.clk(clk_clk),
	.d(sr_21),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_21),
	.prn(vcc));
defparam \jdo[21] .is_wysiwyg = "true";
defparam \jdo[21] .power_up = "low";

dffeas \jdo[20] (
	.clk(clk_clk),
	.d(sr_20),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_20),
	.prn(vcc));
defparam \jdo[20] .is_wysiwyg = "true";
defparam \jdo[20] .power_up = "low";

dffeas \jdo[0] (
	.clk(clk_clk),
	.d(sr_0),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_0),
	.prn(vcc));
defparam \jdo[0] .is_wysiwyg = "true";
defparam \jdo[0] .power_up = "low";

dffeas \jdo[36] (
	.clk(clk_clk),
	.d(sr_36),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_36),
	.prn(vcc));
defparam \jdo[36] .is_wysiwyg = "true";
defparam \jdo[36] .power_up = "low";

dffeas \jdo[37] (
	.clk(clk_clk),
	.d(sr_37),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_37),
	.prn(vcc));
defparam \jdo[37] .is_wysiwyg = "true";
defparam \jdo[37] .power_up = "low";

dffeas \jdo[3] (
	.clk(clk_clk),
	.d(sr_3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_3),
	.prn(vcc));
defparam \jdo[3] .is_wysiwyg = "true";
defparam \jdo[3] .power_up = "low";

dffeas \jdo[19] (
	.clk(clk_clk),
	.d(sr_19),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_19),
	.prn(vcc));
defparam \jdo[19] .is_wysiwyg = "true";
defparam \jdo[19] .power_up = "low";

dffeas \jdo[18] (
	.clk(clk_clk),
	.d(sr_18),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_18),
	.prn(vcc));
defparam \jdo[18] .is_wysiwyg = "true";
defparam \jdo[18] .power_up = "low";

dffeas \jdo[17] (
	.clk(clk_clk),
	.d(sr_17),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_17),
	.prn(vcc));
defparam \jdo[17] .is_wysiwyg = "true";
defparam \jdo[17] .power_up = "low";

dffeas \jdo[25] (
	.clk(clk_clk),
	.d(sr_25),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_25),
	.prn(vcc));
defparam \jdo[25] .is_wysiwyg = "true";
defparam \jdo[25] .power_up = "low";

dffeas \jdo[1] (
	.clk(clk_clk),
	.d(sr_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_1),
	.prn(vcc));
defparam \jdo[1] .is_wysiwyg = "true";
defparam \jdo[1] .power_up = "low";

dffeas \jdo[4] (
	.clk(clk_clk),
	.d(sr_4),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_4),
	.prn(vcc));
defparam \jdo[4] .is_wysiwyg = "true";
defparam \jdo[4] .power_up = "low";

dffeas \jdo[26] (
	.clk(clk_clk),
	.d(sr_26),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_26),
	.prn(vcc));
defparam \jdo[26] .is_wysiwyg = "true";
defparam \jdo[26] .power_up = "low";

dffeas \jdo[27] (
	.clk(clk_clk),
	.d(sr_27),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_27),
	.prn(vcc));
defparam \jdo[27] .is_wysiwyg = "true";
defparam \jdo[27] .power_up = "low";

dffeas \jdo[28] (
	.clk(clk_clk),
	.d(sr_28),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_28),
	.prn(vcc));
defparam \jdo[28] .is_wysiwyg = "true";
defparam \jdo[28] .power_up = "low";

dffeas \jdo[2] (
	.clk(clk_clk),
	.d(sr_2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_2),
	.prn(vcc));
defparam \jdo[2] .is_wysiwyg = "true";
defparam \jdo[2] .power_up = "low";

dffeas \jdo[5] (
	.clk(clk_clk),
	.d(sr_5),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_5),
	.prn(vcc));
defparam \jdo[5] .is_wysiwyg = "true";
defparam \jdo[5] .power_up = "low";

dffeas \jdo[29] (
	.clk(clk_clk),
	.d(sr_29),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_29),
	.prn(vcc));
defparam \jdo[29] .is_wysiwyg = "true";
defparam \jdo[29] .power_up = "low";

dffeas \jdo[30] (
	.clk(clk_clk),
	.d(sr_30),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_30),
	.prn(vcc));
defparam \jdo[30] .is_wysiwyg = "true";
defparam \jdo[30] .power_up = "low";

dffeas \jdo[31] (
	.clk(clk_clk),
	.d(sr_31),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_31),
	.prn(vcc));
defparam \jdo[31] .is_wysiwyg = "true";
defparam \jdo[31] .power_up = "low";

dffeas \jdo[32] (
	.clk(clk_clk),
	.d(sr_32),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_32),
	.prn(vcc));
defparam \jdo[32] .is_wysiwyg = "true";
defparam \jdo[32] .power_up = "low";

dffeas \jdo[33] (
	.clk(clk_clk),
	.d(sr_33),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_33),
	.prn(vcc));
defparam \jdo[33] .is_wysiwyg = "true";
defparam \jdo[33] .power_up = "low";

dffeas \jdo[23] (
	.clk(clk_clk),
	.d(sr_23),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_23),
	.prn(vcc));
defparam \jdo[23] .is_wysiwyg = "true";
defparam \jdo[23] .power_up = "low";

dffeas \jdo[22] (
	.clk(clk_clk),
	.d(sr_22),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_22),
	.prn(vcc));
defparam \jdo[22] .is_wysiwyg = "true";
defparam \jdo[22] .power_up = "low";

dffeas \jdo[6] (
	.clk(clk_clk),
	.d(sr_6),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_6),
	.prn(vcc));
defparam \jdo[6] .is_wysiwyg = "true";
defparam \jdo[6] .power_up = "low";

dffeas \jdo[24] (
	.clk(clk_clk),
	.d(sr_24),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_24),
	.prn(vcc));
defparam \jdo[24] .is_wysiwyg = "true";
defparam \jdo[24] .power_up = "low";

dffeas \jdo[16] (
	.clk(clk_clk),
	.d(sr_16),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_16),
	.prn(vcc));
defparam \jdo[16] .is_wysiwyg = "true";
defparam \jdo[16] .power_up = "low";

dffeas \jdo[7] (
	.clk(clk_clk),
	.d(sr_7),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_7),
	.prn(vcc));
defparam \jdo[7] .is_wysiwyg = "true";
defparam \jdo[7] .power_up = "low";

dffeas \jdo[8] (
	.clk(clk_clk),
	.d(sr_8),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_8),
	.prn(vcc));
defparam \jdo[8] .is_wysiwyg = "true";
defparam \jdo[8] .power_up = "low";

dffeas \jdo[9] (
	.clk(clk_clk),
	.d(sr_9),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_9),
	.prn(vcc));
defparam \jdo[9] .is_wysiwyg = "true";
defparam \jdo[9] .power_up = "low";

dffeas \jdo[10] (
	.clk(clk_clk),
	.d(sr_10),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_10),
	.prn(vcc));
defparam \jdo[10] .is_wysiwyg = "true";
defparam \jdo[10] .power_up = "low";

dffeas \jdo[14] (
	.clk(clk_clk),
	.d(sr_14),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_14),
	.prn(vcc));
defparam \jdo[14] .is_wysiwyg = "true";
defparam \jdo[14] .power_up = "low";

dffeas \jdo[13] (
	.clk(clk_clk),
	.d(sr_13),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_13),
	.prn(vcc));
defparam \jdo[13] .is_wysiwyg = "true";
defparam \jdo[13] .power_up = "low";

dffeas \jdo[11] (
	.clk(clk_clk),
	.d(sr_11),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_11),
	.prn(vcc));
defparam \jdo[11] .is_wysiwyg = "true";
defparam \jdo[11] .power_up = "low";

dffeas \jdo[12] (
	.clk(clk_clk),
	.d(sr_12),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_12),
	.prn(vcc));
defparam \jdo[12] .is_wysiwyg = "true";
defparam \jdo[12] .power_up = "low";

dffeas \jdo[15] (
	.clk(clk_clk),
	.d(sr_15),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_15),
	.prn(vcc));
defparam \jdo[15] .is_wysiwyg = "true";
defparam \jdo[15] .power_up = "low";

dffeas sync2_udr(
	.clk(clk_clk),
	.d(\the_altera_std_synchronizer3|dreg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sync2_udr~q ),
	.prn(vcc));
defparam sync2_udr.is_wysiwyg = "true";
defparam sync2_udr.power_up = "low";

cyclonev_lcell_comb \update_jdo_strobe~0 (
	.dataa(!\sync2_udr~q ),
	.datab(!\the_altera_std_synchronizer3|dreg[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\update_jdo_strobe~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \update_jdo_strobe~0 .extended_lut = "off";
defparam \update_jdo_strobe~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \update_jdo_strobe~0 .shared_arith = "off";

dffeas update_jdo_strobe(
	.clk(clk_clk),
	.d(\update_jdo_strobe~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\update_jdo_strobe~q ),
	.prn(vcc));
defparam update_jdo_strobe.is_wysiwyg = "true";
defparam update_jdo_strobe.power_up = "low";

dffeas sync2_uir(
	.clk(clk_clk),
	.d(\the_altera_std_synchronizer4|dreg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sync2_uir~q ),
	.prn(vcc));
defparam sync2_uir.is_wysiwyg = "true";
defparam sync2_uir.power_up = "low";

cyclonev_lcell_comb \jxuir~0 (
	.dataa(!\sync2_uir~q ),
	.datab(!\the_altera_std_synchronizer4|dreg[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\jxuir~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \jxuir~0 .extended_lut = "off";
defparam \jxuir~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \jxuir~0 .shared_arith = "off";

dffeas jxuir(
	.clk(clk_clk),
	.d(\jxuir~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jxuir~q ),
	.prn(vcc));
defparam jxuir.is_wysiwyg = "true";
defparam jxuir.power_up = "low";

endmodule

module first_nios2_system_altera_std_synchronizer (
	dreg_0,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_0;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module first_nios2_system_altera_std_synchronizer_1 (
	din,
	dreg_0,
	clk)/* synthesis synthesis_greybox=1 */;
input 	din;
output 	dreg_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module first_nios2_system_first_nios2_system_cpu_cpu_debug_slave_tck (
	sr_1,
	sr_2,
	break_readreg_0,
	sr_3,
	break_readreg_1,
	sr_21,
	sr_20,
	sr_4,
	break_readreg_2,
	MonDReg_2,
	sr_22,
	break_readreg_20,
	MonDReg_20,
	break_readreg_19,
	MonDReg_19,
	sr_19,
	sr_18,
	sr_17,
	sr_25,
	sr_5,
	break_readreg_3,
	sr_26,
	sr_27,
	sr_28,
	sr_23,
	break_readreg_21,
	MonDReg_21,
	break_readreg_18,
	break_readreg_17,
	MonDReg_17,
	break_readreg_16,
	MonDReg_16,
	break_readreg_24,
	MonDReg_24,
	sr_6,
	break_readreg_4,
	break_readreg_25,
	MonDReg_25,
	break_readreg_26,
	MonDReg_26,
	sr_29,
	break_readreg_27,
	MonDReg_27,
	sr_30,
	sr_32,
	sr_24,
	break_readreg_22,
	break_readreg_5,
	break_readreg_28,
	MonDReg_28,
	break_readreg_29,
	MonDReg_30,
	break_readreg_30,
	break_readreg_31,
	MonDReg_31,
	break_readreg_23,
	MonDReg_23,
	sr_16,
	MonDReg_6,
	MonDReg_7,
	sr_8,
	break_readreg_6,
	MonDReg_11,
	MonDReg_10,
	MonDReg_9,
	MonDReg_13,
	MonDReg_14,
	break_readreg_15,
	sr_9,
	break_readreg_7,
	sr_10,
	break_readreg_8,
	sr_14,
	sr_13,
	sr_11,
	sr_12,
	break_readreg_9,
	break_readreg_13,
	break_readreg_12,
	break_readreg_10,
	break_readreg_11,
	break_readreg_14,
	sr_0,
	ir_out_0,
	ir_out_1,
	virtual_state_sdr,
	W_debug_mode,
	MonDReg_0,
	virtual_state_uir,
	monitor_ready,
	MonDReg_1,
	sr_34,
	sr_35,
	sr_36,
	sr_37,
	monitor_error,
	virtual_state_cdr,
	MonDReg_3,
	MonDReg_18,
	MonDReg_4,
	sr_31,
	sr_33,
	MonDReg_22,
	sr_7,
	MonDReg_5,
	MonDReg_29,
	resetlatch,
	MonDReg_8,
	MonDReg_15,
	MonDReg_12,
	sr_15,
	altera_internal_jtag,
	altera_internal_jtag1,
	state_4,
	virtual_ir_scan_reg,
	state_3,
	splitter_nodes_receive_1_3,
	irf_reg_0_2,
	irf_reg_1_2)/* synthesis synthesis_greybox=1 */;
output 	sr_1;
output 	sr_2;
input 	break_readreg_0;
output 	sr_3;
input 	break_readreg_1;
output 	sr_21;
output 	sr_20;
output 	sr_4;
input 	break_readreg_2;
input 	MonDReg_2;
output 	sr_22;
input 	break_readreg_20;
input 	MonDReg_20;
input 	break_readreg_19;
input 	MonDReg_19;
output 	sr_19;
output 	sr_18;
output 	sr_17;
output 	sr_25;
output 	sr_5;
input 	break_readreg_3;
output 	sr_26;
output 	sr_27;
output 	sr_28;
output 	sr_23;
input 	break_readreg_21;
input 	MonDReg_21;
input 	break_readreg_18;
input 	break_readreg_17;
input 	MonDReg_17;
input 	break_readreg_16;
input 	MonDReg_16;
input 	break_readreg_24;
input 	MonDReg_24;
output 	sr_6;
input 	break_readreg_4;
input 	break_readreg_25;
input 	MonDReg_25;
input 	break_readreg_26;
input 	MonDReg_26;
output 	sr_29;
input 	break_readreg_27;
input 	MonDReg_27;
output 	sr_30;
output 	sr_32;
output 	sr_24;
input 	break_readreg_22;
input 	break_readreg_5;
input 	break_readreg_28;
input 	MonDReg_28;
input 	break_readreg_29;
input 	MonDReg_30;
input 	break_readreg_30;
input 	break_readreg_31;
input 	MonDReg_31;
input 	break_readreg_23;
input 	MonDReg_23;
output 	sr_16;
input 	MonDReg_6;
input 	MonDReg_7;
output 	sr_8;
input 	break_readreg_6;
input 	MonDReg_11;
input 	MonDReg_10;
input 	MonDReg_9;
input 	MonDReg_13;
input 	MonDReg_14;
input 	break_readreg_15;
output 	sr_9;
input 	break_readreg_7;
output 	sr_10;
input 	break_readreg_8;
output 	sr_14;
output 	sr_13;
output 	sr_11;
output 	sr_12;
input 	break_readreg_9;
input 	break_readreg_13;
input 	break_readreg_12;
input 	break_readreg_10;
input 	break_readreg_11;
input 	break_readreg_14;
output 	sr_0;
output 	ir_out_0;
output 	ir_out_1;
input 	virtual_state_sdr;
input 	W_debug_mode;
input 	MonDReg_0;
input 	virtual_state_uir;
input 	monitor_ready;
input 	MonDReg_1;
output 	sr_34;
output 	sr_35;
output 	sr_36;
output 	sr_37;
input 	monitor_error;
input 	virtual_state_cdr;
input 	MonDReg_3;
input 	MonDReg_18;
input 	MonDReg_4;
output 	sr_31;
output 	sr_33;
input 	MonDReg_22;
output 	sr_7;
input 	MonDReg_5;
input 	MonDReg_29;
input 	resetlatch;
input 	MonDReg_8;
input 	MonDReg_15;
input 	MonDReg_12;
output 	sr_15;
input 	altera_internal_jtag;
input 	altera_internal_jtag1;
input 	state_4;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	splitter_nodes_receive_1_3;
input 	irf_reg_0_2;
input 	irf_reg_1_2;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \the_altera_std_synchronizer2|dreg[0]~q ;
wire \the_altera_std_synchronizer1|dreg[0]~q ;
wire \sr~8_combout ;
wire \sr[1]~9_combout ;
wire \sr[1]~10_combout ;
wire \sr~11_combout ;
wire \sr~12_combout ;
wire \sr~16_combout ;
wire \sr[29]~17_combout ;
wire \sr[29]~14_combout ;
wire \sr~18_combout ;
wire \sr~19_combout ;
wire \sr~23_combout ;
wire \sr~24_combout ;
wire \sr~25_combout ;
wire \sr~26_combout ;
wire \sr~27_combout ;
wire \sr~28_combout ;
wire \sr~29_combout ;
wire \sr~30_combout ;
wire \sr~31_combout ;
wire \sr~32_combout ;
wire \sr~33_combout ;
wire \sr~34_combout ;
wire \sr~35_combout ;
wire \sr~40_combout ;
wire \sr~42_combout ;
wire \sr~45_combout ;
wire \sr~46_combout ;
wire \sr~47_combout ;
wire \sr~48_combout ;
wire \sr~49_combout ;
wire \sr~50_combout ;
wire \sr~51_combout ;
wire \sr~52_combout ;
wire \sr~5_combout ;
wire \sr~6_combout ;
wire \DRsize.000~q ;
wire \sr~7_combout ;
wire \Mux37~0_combout ;
wire \sr~13_combout ;
wire \DRsize.100~q ;
wire \sr~56_combout ;
wire \sr~15_combout ;
wire \sr~20_combout ;
wire \sr[37]~21_combout ;
wire \sr~22_combout ;
wire \sr[29]~36_combout ;
wire \sr~37_combout ;
wire \sr~38_combout ;
wire \sr~39_combout ;
wire \sr~41_combout ;
wire \sr~43_combout ;
wire \sr~44_combout ;
wire \sr[29]~55_combout ;
wire \DRsize.010~q ;
wire \sr~53_combout ;
wire \sr~54_combout ;


first_nios2_system_altera_std_synchronizer_3 the_altera_std_synchronizer2(
	.dreg_0(\the_altera_std_synchronizer2|dreg[0]~q ),
	.din(monitor_ready),
	.clk(altera_internal_jtag));

first_nios2_system_altera_std_synchronizer_2 the_altera_std_synchronizer1(
	.dreg_0(\the_altera_std_synchronizer1|dreg[0]~q ),
	.din(W_debug_mode),
	.clk(altera_internal_jtag));

dffeas \sr[1] (
	.clk(altera_internal_jtag),
	.d(\sr~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[1]~9_combout ),
	.sload(gnd),
	.ena(\sr[1]~10_combout ),
	.q(sr_1),
	.prn(vcc));
defparam \sr[1] .is_wysiwyg = "true";
defparam \sr[1] .power_up = "low";

dffeas \sr[2] (
	.clk(altera_internal_jtag),
	.d(\sr~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[1]~9_combout ),
	.sload(gnd),
	.ena(\sr[1]~10_combout ),
	.q(sr_2),
	.prn(vcc));
defparam \sr[2] .is_wysiwyg = "true";
defparam \sr[2] .power_up = "low";

dffeas \sr[3] (
	.clk(altera_internal_jtag),
	.d(\sr~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[1]~9_combout ),
	.sload(gnd),
	.ena(\sr[1]~10_combout ),
	.q(sr_3),
	.prn(vcc));
defparam \sr[3] .is_wysiwyg = "true";
defparam \sr[3] .power_up = "low";

dffeas \sr[21] (
	.clk(altera_internal_jtag),
	.d(\sr~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[29]~17_combout ),
	.sload(gnd),
	.ena(\sr[29]~14_combout ),
	.q(sr_21),
	.prn(vcc));
defparam \sr[21] .is_wysiwyg = "true";
defparam \sr[21] .power_up = "low";

dffeas \sr[20] (
	.clk(altera_internal_jtag),
	.d(\sr~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[29]~17_combout ),
	.sload(gnd),
	.ena(\sr[29]~14_combout ),
	.q(sr_20),
	.prn(vcc));
defparam \sr[20] .is_wysiwyg = "true";
defparam \sr[20] .power_up = "low";

dffeas \sr[4] (
	.clk(altera_internal_jtag),
	.d(\sr~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[1]~9_combout ),
	.sload(gnd),
	.ena(\sr[1]~10_combout ),
	.q(sr_4),
	.prn(vcc));
defparam \sr[4] .is_wysiwyg = "true";
defparam \sr[4] .power_up = "low";

dffeas \sr[22] (
	.clk(altera_internal_jtag),
	.d(\sr~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[29]~17_combout ),
	.sload(gnd),
	.ena(\sr[29]~14_combout ),
	.q(sr_22),
	.prn(vcc));
defparam \sr[22] .is_wysiwyg = "true";
defparam \sr[22] .power_up = "low";

dffeas \sr[19] (
	.clk(altera_internal_jtag),
	.d(\sr~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[29]~17_combout ),
	.sload(gnd),
	.ena(\sr[29]~14_combout ),
	.q(sr_19),
	.prn(vcc));
defparam \sr[19] .is_wysiwyg = "true";
defparam \sr[19] .power_up = "low";

dffeas \sr[18] (
	.clk(altera_internal_jtag),
	.d(\sr~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[29]~17_combout ),
	.sload(gnd),
	.ena(\sr[29]~14_combout ),
	.q(sr_18),
	.prn(vcc));
defparam \sr[18] .is_wysiwyg = "true";
defparam \sr[18] .power_up = "low";

dffeas \sr[17] (
	.clk(altera_internal_jtag),
	.d(\sr~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[29]~17_combout ),
	.sload(gnd),
	.ena(\sr[29]~14_combout ),
	.q(sr_17),
	.prn(vcc));
defparam \sr[17] .is_wysiwyg = "true";
defparam \sr[17] .power_up = "low";

dffeas \sr[25] (
	.clk(altera_internal_jtag),
	.d(\sr~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[29]~17_combout ),
	.sload(gnd),
	.ena(\sr[29]~14_combout ),
	.q(sr_25),
	.prn(vcc));
defparam \sr[25] .is_wysiwyg = "true";
defparam \sr[25] .power_up = "low";

dffeas \sr[5] (
	.clk(altera_internal_jtag),
	.d(\sr~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[1]~9_combout ),
	.sload(gnd),
	.ena(\sr[1]~10_combout ),
	.q(sr_5),
	.prn(vcc));
defparam \sr[5] .is_wysiwyg = "true";
defparam \sr[5] .power_up = "low";

dffeas \sr[26] (
	.clk(altera_internal_jtag),
	.d(\sr~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[29]~17_combout ),
	.sload(gnd),
	.ena(\sr[29]~14_combout ),
	.q(sr_26),
	.prn(vcc));
defparam \sr[26] .is_wysiwyg = "true";
defparam \sr[26] .power_up = "low";

dffeas \sr[27] (
	.clk(altera_internal_jtag),
	.d(\sr~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[29]~17_combout ),
	.sload(gnd),
	.ena(\sr[29]~14_combout ),
	.q(sr_27),
	.prn(vcc));
defparam \sr[27] .is_wysiwyg = "true";
defparam \sr[27] .power_up = "low";

dffeas \sr[28] (
	.clk(altera_internal_jtag),
	.d(\sr~31_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[29]~17_combout ),
	.sload(gnd),
	.ena(\sr[29]~14_combout ),
	.q(sr_28),
	.prn(vcc));
defparam \sr[28] .is_wysiwyg = "true";
defparam \sr[28] .power_up = "low";

dffeas \sr[23] (
	.clk(altera_internal_jtag),
	.d(\sr~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[29]~17_combout ),
	.sload(gnd),
	.ena(\sr[29]~14_combout ),
	.q(sr_23),
	.prn(vcc));
defparam \sr[23] .is_wysiwyg = "true";
defparam \sr[23] .power_up = "low";

dffeas \sr[6] (
	.clk(altera_internal_jtag),
	.d(\sr~33_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[1]~9_combout ),
	.sload(gnd),
	.ena(\sr[1]~10_combout ),
	.q(sr_6),
	.prn(vcc));
defparam \sr[6] .is_wysiwyg = "true";
defparam \sr[6] .power_up = "low";

dffeas \sr[29] (
	.clk(altera_internal_jtag),
	.d(\sr~34_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[29]~17_combout ),
	.sload(gnd),
	.ena(\sr[29]~14_combout ),
	.q(sr_29),
	.prn(vcc));
defparam \sr[29] .is_wysiwyg = "true";
defparam \sr[29] .power_up = "low";

dffeas \sr[30] (
	.clk(altera_internal_jtag),
	.d(\sr~35_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[29]~17_combout ),
	.sload(gnd),
	.ena(\sr[29]~14_combout ),
	.q(sr_30),
	.prn(vcc));
defparam \sr[30] .is_wysiwyg = "true";
defparam \sr[30] .power_up = "low";

dffeas \sr[32] (
	.clk(altera_internal_jtag),
	.d(\sr~40_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[29]~17_combout ),
	.sload(gnd),
	.ena(\sr[29]~14_combout ),
	.q(sr_32),
	.prn(vcc));
defparam \sr[32] .is_wysiwyg = "true";
defparam \sr[32] .power_up = "low";

dffeas \sr[24] (
	.clk(altera_internal_jtag),
	.d(\sr~42_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[29]~17_combout ),
	.sload(gnd),
	.ena(\sr[29]~14_combout ),
	.q(sr_24),
	.prn(vcc));
defparam \sr[24] .is_wysiwyg = "true";
defparam \sr[24] .power_up = "low";

dffeas \sr[16] (
	.clk(altera_internal_jtag),
	.d(\sr~45_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[29]~17_combout ),
	.sload(gnd),
	.ena(\sr[29]~14_combout ),
	.q(sr_16),
	.prn(vcc));
defparam \sr[16] .is_wysiwyg = "true";
defparam \sr[16] .power_up = "low";

dffeas \sr[8] (
	.clk(altera_internal_jtag),
	.d(\sr~46_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[1]~9_combout ),
	.sload(gnd),
	.ena(\sr[1]~10_combout ),
	.q(sr_8),
	.prn(vcc));
defparam \sr[8] .is_wysiwyg = "true";
defparam \sr[8] .power_up = "low";

dffeas \sr[9] (
	.clk(altera_internal_jtag),
	.d(\sr~47_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[1]~9_combout ),
	.sload(gnd),
	.ena(\sr[1]~10_combout ),
	.q(sr_9),
	.prn(vcc));
defparam \sr[9] .is_wysiwyg = "true";
defparam \sr[9] .power_up = "low";

dffeas \sr[10] (
	.clk(altera_internal_jtag),
	.d(\sr~48_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[1]~9_combout ),
	.sload(gnd),
	.ena(\sr[1]~10_combout ),
	.q(sr_10),
	.prn(vcc));
defparam \sr[10] .is_wysiwyg = "true";
defparam \sr[10] .power_up = "low";

dffeas \sr[14] (
	.clk(altera_internal_jtag),
	.d(\sr~49_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[1]~9_combout ),
	.sload(gnd),
	.ena(\sr[1]~10_combout ),
	.q(sr_14),
	.prn(vcc));
defparam \sr[14] .is_wysiwyg = "true";
defparam \sr[14] .power_up = "low";

dffeas \sr[13] (
	.clk(altera_internal_jtag),
	.d(\sr~50_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[1]~9_combout ),
	.sload(gnd),
	.ena(\sr[1]~10_combout ),
	.q(sr_13),
	.prn(vcc));
defparam \sr[13] .is_wysiwyg = "true";
defparam \sr[13] .power_up = "low";

dffeas \sr[11] (
	.clk(altera_internal_jtag),
	.d(\sr~51_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[1]~9_combout ),
	.sload(gnd),
	.ena(\sr[1]~10_combout ),
	.q(sr_11),
	.prn(vcc));
defparam \sr[11] .is_wysiwyg = "true";
defparam \sr[11] .power_up = "low";

dffeas \sr[12] (
	.clk(altera_internal_jtag),
	.d(\sr~52_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[1]~9_combout ),
	.sload(gnd),
	.ena(\sr[1]~10_combout ),
	.q(sr_12),
	.prn(vcc));
defparam \sr[12] .is_wysiwyg = "true";
defparam \sr[12] .power_up = "low";

dffeas \sr[0] (
	.clk(altera_internal_jtag),
	.d(\sr~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(sr_0),
	.prn(vcc));
defparam \sr[0] .is_wysiwyg = "true";
defparam \sr[0] .power_up = "low";

dffeas \ir_out[0] (
	.clk(altera_internal_jtag),
	.d(\the_altera_std_synchronizer2|dreg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ir_out_0),
	.prn(vcc));
defparam \ir_out[0] .is_wysiwyg = "true";
defparam \ir_out[0] .power_up = "low";

dffeas \ir_out[1] (
	.clk(altera_internal_jtag),
	.d(\the_altera_std_synchronizer1|dreg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ir_out_1),
	.prn(vcc));
defparam \ir_out[1] .is_wysiwyg = "true";
defparam \ir_out[1] .power_up = "low";

dffeas \sr[34] (
	.clk(altera_internal_jtag),
	.d(\sr~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[29]~14_combout ),
	.q(sr_34),
	.prn(vcc));
defparam \sr[34] .is_wysiwyg = "true";
defparam \sr[34] .power_up = "low";

dffeas \sr[35] (
	.clk(altera_internal_jtag),
	.d(\sr~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(sr_35),
	.prn(vcc));
defparam \sr[35] .is_wysiwyg = "true";
defparam \sr[35] .power_up = "low";

dffeas \sr[36] (
	.clk(altera_internal_jtag),
	.d(\sr~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[37]~21_combout ),
	.q(sr_36),
	.prn(vcc));
defparam \sr[36] .is_wysiwyg = "true";
defparam \sr[36] .power_up = "low";

dffeas \sr[37] (
	.clk(altera_internal_jtag),
	.d(\sr~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[37]~21_combout ),
	.q(sr_37),
	.prn(vcc));
defparam \sr[37] .is_wysiwyg = "true";
defparam \sr[37] .power_up = "low";

dffeas \sr[31] (
	.clk(altera_internal_jtag),
	.d(\sr~39_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(sr_31),
	.prn(vcc));
defparam \sr[31] .is_wysiwyg = "true";
defparam \sr[31] .power_up = "low";

dffeas \sr[33] (
	.clk(altera_internal_jtag),
	.d(\sr~41_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[29]~14_combout ),
	.q(sr_33),
	.prn(vcc));
defparam \sr[33] .is_wysiwyg = "true";
defparam \sr[33] .power_up = "low";

dffeas \sr[7] (
	.clk(altera_internal_jtag),
	.d(\sr~44_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(sr_7),
	.prn(vcc));
defparam \sr[7] .is_wysiwyg = "true";
defparam \sr[7] .power_up = "low";

dffeas \sr[15] (
	.clk(altera_internal_jtag),
	.d(\sr~54_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(sr_15),
	.prn(vcc));
defparam \sr[15] .is_wysiwyg = "true";
defparam \sr[15] .power_up = "low";

cyclonev_lcell_comb \sr~8 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_2),
	.datad(!break_readreg_0),
	.datae(!MonDReg_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~8 .extended_lut = "off";
defparam \sr~8 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~8 .shared_arith = "off";

cyclonev_lcell_comb \sr[1]~9 (
	.dataa(!state_4),
	.datab(!virtual_ir_scan_reg),
	.datac(!splitter_nodes_receive_1_3),
	.datad(!irf_reg_0_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr[1]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr[1]~9 .extended_lut = "off";
defparam \sr[1]~9 .lut_mask = 64'hFBFFFBFFFBFFFBFF;
defparam \sr[1]~9 .shared_arith = "off";

cyclonev_lcell_comb \sr[1]~10 (
	.dataa(!state_4),
	.datab(!virtual_ir_scan_reg),
	.datac(!splitter_nodes_receive_1_3),
	.datad(!state_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr[1]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr[1]~10 .extended_lut = "off";
defparam \sr[1]~10 .lut_mask = 64'hDFFFDFFFDFFFDFFF;
defparam \sr[1]~10 .shared_arith = "off";

cyclonev_lcell_comb \sr~11 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_3),
	.datad(!break_readreg_1),
	.datae(!MonDReg_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~11 .extended_lut = "off";
defparam \sr~11 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~11 .shared_arith = "off";

cyclonev_lcell_comb \sr~12 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_4),
	.datad(!break_readreg_2),
	.datae(!MonDReg_2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~12 .extended_lut = "off";
defparam \sr~12 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~12 .shared_arith = "off";

cyclonev_lcell_comb \sr~16 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_22),
	.datad(!break_readreg_20),
	.datae(!MonDReg_20),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~16 .extended_lut = "off";
defparam \sr~16 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~16 .shared_arith = "off";

cyclonev_lcell_comb \sr[29]~17 (
	.dataa(!state_4),
	.datab(!virtual_ir_scan_reg),
	.datac(!splitter_nodes_receive_1_3),
	.datad(!irf_reg_0_2),
	.datae(!irf_reg_1_2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr[29]~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr[29]~17 .extended_lut = "off";
defparam \sr[29]~17 .lut_mask = 64'hFFFFFBFFFFFFFBFF;
defparam \sr[29]~17 .shared_arith = "off";

cyclonev_lcell_comb \sr[29]~14 (
	.dataa(!state_4),
	.datab(!virtual_ir_scan_reg),
	.datac(!splitter_nodes_receive_1_3),
	.datad(!state_3),
	.datae(!irf_reg_0_2),
	.dataf(!irf_reg_1_2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr[29]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr[29]~14 .extended_lut = "off";
defparam \sr[29]~14 .lut_mask = 64'hFFFFFFFFFFFFDFFF;
defparam \sr[29]~14 .shared_arith = "off";

cyclonev_lcell_comb \sr~18 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_21),
	.datad(!break_readreg_19),
	.datae(!MonDReg_19),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~18 .extended_lut = "off";
defparam \sr~18 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~18 .shared_arith = "off";

cyclonev_lcell_comb \sr~19 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_5),
	.datad(!break_readreg_3),
	.datae(!MonDReg_3),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~19 .extended_lut = "off";
defparam \sr~19 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~19 .shared_arith = "off";

cyclonev_lcell_comb \sr~23 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_23),
	.datad(!break_readreg_21),
	.datae(!MonDReg_21),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~23 .extended_lut = "off";
defparam \sr~23 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~23 .shared_arith = "off";

cyclonev_lcell_comb \sr~24 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_20),
	.datad(!break_readreg_18),
	.datae(!MonDReg_18),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~24 .extended_lut = "off";
defparam \sr~24 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~24 .shared_arith = "off";

cyclonev_lcell_comb \sr~25 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_19),
	.datad(!break_readreg_17),
	.datae(!MonDReg_17),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~25 .extended_lut = "off";
defparam \sr~25 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~25 .shared_arith = "off";

cyclonev_lcell_comb \sr~26 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_18),
	.datad(!break_readreg_16),
	.datae(!MonDReg_16),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~26 .extended_lut = "off";
defparam \sr~26 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~26 .shared_arith = "off";

cyclonev_lcell_comb \sr~27 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_26),
	.datad(!break_readreg_24),
	.datae(!MonDReg_24),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~27 .extended_lut = "off";
defparam \sr~27 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~27 .shared_arith = "off";

cyclonev_lcell_comb \sr~28 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_6),
	.datad(!break_readreg_4),
	.datae(!MonDReg_4),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~28 .extended_lut = "off";
defparam \sr~28 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~28 .shared_arith = "off";

cyclonev_lcell_comb \sr~29 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_27),
	.datad(!break_readreg_25),
	.datae(!MonDReg_25),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~29 .extended_lut = "off";
defparam \sr~29 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~29 .shared_arith = "off";

cyclonev_lcell_comb \sr~30 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_28),
	.datad(!break_readreg_26),
	.datae(!MonDReg_26),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~30 .extended_lut = "off";
defparam \sr~30 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~30 .shared_arith = "off";

cyclonev_lcell_comb \sr~31 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_29),
	.datad(!break_readreg_27),
	.datae(!MonDReg_27),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~31 .extended_lut = "off";
defparam \sr~31 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~31 .shared_arith = "off";

cyclonev_lcell_comb \sr~32 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_24),
	.datad(!break_readreg_22),
	.datae(!MonDReg_22),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~32_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~32 .extended_lut = "off";
defparam \sr~32 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~32 .shared_arith = "off";

cyclonev_lcell_comb \sr~33 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_7),
	.datad(!break_readreg_5),
	.datae(!MonDReg_5),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~33_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~33 .extended_lut = "off";
defparam \sr~33 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~33 .shared_arith = "off";

cyclonev_lcell_comb \sr~34 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_30),
	.datad(!break_readreg_28),
	.datae(!MonDReg_28),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~34_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~34 .extended_lut = "off";
defparam \sr~34 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~34 .shared_arith = "off";

cyclonev_lcell_comb \sr~35 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_31),
	.datad(!break_readreg_29),
	.datae(!MonDReg_29),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~35_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~35 .extended_lut = "off";
defparam \sr~35 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~35 .shared_arith = "off";

cyclonev_lcell_comb \sr~40 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_33),
	.datad(!break_readreg_31),
	.datae(!MonDReg_31),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~40_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~40 .extended_lut = "off";
defparam \sr~40 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~40 .shared_arith = "off";

cyclonev_lcell_comb \sr~42 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_25),
	.datad(!break_readreg_23),
	.datae(!MonDReg_23),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~42_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~42 .extended_lut = "off";
defparam \sr~42 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~42 .shared_arith = "off";

cyclonev_lcell_comb \sr~45 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_17),
	.datad(!MonDReg_15),
	.datae(!break_readreg_15),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~45_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~45 .extended_lut = "off";
defparam \sr~45 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~45 .shared_arith = "off";

cyclonev_lcell_comb \sr~46 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!MonDReg_7),
	.datad(!sr_9),
	.datae(!break_readreg_7),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~46_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~46 .extended_lut = "off";
defparam \sr~46 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~46 .shared_arith = "off";

cyclonev_lcell_comb \sr~47 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!MonDReg_8),
	.datad(!sr_10),
	.datae(!break_readreg_8),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~47_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~47 .extended_lut = "off";
defparam \sr~47 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~47 .shared_arith = "off";

cyclonev_lcell_comb \sr~48 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!MonDReg_9),
	.datad(!sr_11),
	.datae(!break_readreg_9),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~48_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~48 .extended_lut = "off";
defparam \sr~48 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~48 .shared_arith = "off";

cyclonev_lcell_comb \sr~49 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!MonDReg_13),
	.datad(!sr_15),
	.datae(!break_readreg_13),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~49_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~49 .extended_lut = "off";
defparam \sr~49 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~49 .shared_arith = "off";

cyclonev_lcell_comb \sr~50 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!MonDReg_12),
	.datad(!sr_14),
	.datae(!break_readreg_12),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~50_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~50 .extended_lut = "off";
defparam \sr~50 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~50 .shared_arith = "off";

cyclonev_lcell_comb \sr~51 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!MonDReg_10),
	.datad(!sr_12),
	.datae(!break_readreg_10),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~51_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~51 .extended_lut = "off";
defparam \sr~51 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~51 .shared_arith = "off";

cyclonev_lcell_comb \sr~52 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!MonDReg_11),
	.datad(!sr_13),
	.datae(!break_readreg_11),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~52_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~52 .extended_lut = "off";
defparam \sr~52 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~52 .shared_arith = "off";

cyclonev_lcell_comb \sr~5 (
	.dataa(!sr_0),
	.datab(!virtual_ir_scan_reg),
	.datac(!splitter_nodes_receive_1_3),
	.datad(!state_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~5 .extended_lut = "off";
defparam \sr~5 .lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam \sr~5 .shared_arith = "off";

cyclonev_lcell_comb \sr~6 (
	.dataa(!virtual_ir_scan_reg),
	.datab(!splitter_nodes_receive_1_3),
	.datac(!state_3),
	.datad(!\the_altera_std_synchronizer2|dreg[0]~q ),
	.datae(!irf_reg_0_2),
	.dataf(!irf_reg_1_2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~6 .extended_lut = "off";
defparam \sr~6 .lut_mask = 64'hFFFFFFFFFFFFBFFF;
defparam \sr~6 .shared_arith = "off";

dffeas \DRsize.000 (
	.clk(altera_internal_jtag),
	.d(vcc),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(virtual_state_uir),
	.q(\DRsize.000~q ),
	.prn(vcc));
defparam \DRsize.000 .is_wysiwyg = "true";
defparam \DRsize.000 .power_up = "low";

cyclonev_lcell_comb \sr~7 (
	.dataa(!virtual_state_sdr),
	.datab(!\sr~5_combout ),
	.datac(!\sr~6_combout ),
	.datad(!sr_1),
	.datae(!\DRsize.000~q ),
	.dataf(!altera_internal_jtag1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~7 .extended_lut = "off";
defparam \sr~7 .lut_mask = 64'h7FFFBFFFFFFFFFFF;
defparam \sr~7 .shared_arith = "off";

cyclonev_lcell_comb \Mux37~0 (
	.dataa(!irf_reg_0_2),
	.datab(!irf_reg_1_2),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux37~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux37~0 .extended_lut = "off";
defparam \Mux37~0 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \Mux37~0 .shared_arith = "off";

cyclonev_lcell_comb \sr~13 (
	.dataa(!virtual_state_sdr),
	.datab(!\Mux37~0_combout ),
	.datac(!sr_35),
	.datad(!monitor_error),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~13 .extended_lut = "off";
defparam \sr~13 .lut_mask = 64'h27FF27FF27FF27FF;
defparam \sr~13 .shared_arith = "off";

dffeas \DRsize.100 (
	.clk(altera_internal_jtag),
	.d(\Mux37~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(virtual_state_uir),
	.q(\DRsize.100~q ),
	.prn(vcc));
defparam \DRsize.100 .is_wysiwyg = "true";
defparam \DRsize.100 .power_up = "low";

cyclonev_lcell_comb \sr~56 (
	.dataa(!virtual_state_cdr),
	.datab(!sr_35),
	.datac(!irf_reg_0_2),
	.datad(!irf_reg_1_2),
	.datae(!\the_altera_std_synchronizer1|dreg[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~56_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~56 .extended_lut = "off";
defparam \sr~56 .lut_mask = 64'hB77BFFFFB77BFFFF;
defparam \sr~56 .shared_arith = "off";

cyclonev_lcell_comb \sr~15 (
	.dataa(!virtual_state_sdr),
	.datab(!altera_internal_jtag1),
	.datac(!sr_36),
	.datad(!\DRsize.100~q ),
	.datae(!\sr~56_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~15 .extended_lut = "off";
defparam \sr~15 .lut_mask = 64'h7FBFFFFF7FBFFFFF;
defparam \sr~15 .shared_arith = "off";

cyclonev_lcell_comb \sr~20 (
	.dataa(!state_4),
	.datab(!virtual_ir_scan_reg),
	.datac(!splitter_nodes_receive_1_3),
	.datad(!sr_37),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~20 .extended_lut = "off";
defparam \sr~20 .lut_mask = 64'hDFFFDFFFDFFFDFFF;
defparam \sr~20 .shared_arith = "off";

cyclonev_lcell_comb \sr[37]~21 (
	.dataa(!state_4),
	.datab(!virtual_ir_scan_reg),
	.datac(!splitter_nodes_receive_1_3),
	.datad(!state_3),
	.datae(!irf_reg_0_2),
	.dataf(!irf_reg_1_2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr[37]~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr[37]~21 .extended_lut = "off";
defparam \sr[37]~21 .lut_mask = 64'hDFFFFFFFFFFFDFFF;
defparam \sr[37]~21 .shared_arith = "off";

cyclonev_lcell_comb \sr~22 (
	.dataa(!state_4),
	.datab(!virtual_ir_scan_reg),
	.datac(!splitter_nodes_receive_1_3),
	.datad(!altera_internal_jtag1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~22 .extended_lut = "off";
defparam \sr~22 .lut_mask = 64'hDFFFDFFFDFFFDFFF;
defparam \sr~22 .shared_arith = "off";

cyclonev_lcell_comb \sr[29]~36 (
	.dataa(!virtual_ir_scan_reg),
	.datab(!splitter_nodes_receive_1_3),
	.datac(!state_3),
	.datad(!irf_reg_0_2),
	.datae(!irf_reg_1_2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr[29]~36_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr[29]~36 .extended_lut = "off";
defparam \sr[29]~36 .lut_mask = 64'hFFFFFFBFFFFFFFBF;
defparam \sr[29]~36 .shared_arith = "off";

cyclonev_lcell_comb \sr~37 (
	.dataa(!irf_reg_1_2),
	.datab(!MonDReg_30),
	.datac(!break_readreg_30),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~37_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~37 .extended_lut = "off";
defparam \sr~37 .lut_mask = 64'h2727272727272727;
defparam \sr~37 .shared_arith = "off";

cyclonev_lcell_comb \sr~38 (
	.dataa(!virtual_ir_scan_reg),
	.datab(!splitter_nodes_receive_1_3),
	.datac(!state_3),
	.datad(!irf_reg_0_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~38_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~38 .extended_lut = "off";
defparam \sr~38 .lut_mask = 64'hFFBFFFBFFFBFFFBF;
defparam \sr~38 .shared_arith = "off";

cyclonev_lcell_comb \sr~39 (
	.dataa(!virtual_state_sdr),
	.datab(!\sr[29]~36_combout ),
	.datac(!sr_31),
	.datad(!sr_32),
	.datae(!\sr~37_combout ),
	.dataf(!\sr~38_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~39_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~39 .extended_lut = "off";
defparam \sr~39 .lut_mask = 64'h8DFFFFFFFFFFFFFF;
defparam \sr~39 .shared_arith = "off";

cyclonev_lcell_comb \sr~41 (
	.dataa(!virtual_state_sdr),
	.datab(!\Mux37~0_combout ),
	.datac(!sr_34),
	.datad(!resetlatch),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~41_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~41 .extended_lut = "off";
defparam \sr~41 .lut_mask = 64'h27FF27FF27FF27FF;
defparam \sr~41 .shared_arith = "off";

cyclonev_lcell_comb \sr~43 (
	.dataa(!irf_reg_1_2),
	.datab(!MonDReg_6),
	.datac(!break_readreg_6),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~43_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~43 .extended_lut = "off";
defparam \sr~43 .lut_mask = 64'h2727272727272727;
defparam \sr~43 .shared_arith = "off";

cyclonev_lcell_comb \sr~44 (
	.dataa(!virtual_state_sdr),
	.datab(!virtual_state_cdr),
	.datac(!irf_reg_0_2),
	.datad(!sr_7),
	.datae(!sr_8),
	.dataf(!\sr~43_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~44_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~44 .extended_lut = "off";
defparam \sr~44 .lut_mask = 64'hF6FFFFFFFFFFFFFF;
defparam \sr~44 .shared_arith = "off";

cyclonev_lcell_comb \sr[29]~55 (
	.dataa(!irf_reg_0_2),
	.datab(!irf_reg_1_2),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr[29]~55_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr[29]~55 .extended_lut = "off";
defparam \sr[29]~55 .lut_mask = 64'h7777777777777777;
defparam \sr[29]~55 .shared_arith = "off";

dffeas \DRsize.010 (
	.clk(altera_internal_jtag),
	.d(\sr[29]~55_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(virtual_state_uir),
	.q(\DRsize.010~q ),
	.prn(vcc));
defparam \DRsize.010 .is_wysiwyg = "true";
defparam \DRsize.010 .power_up = "low";

cyclonev_lcell_comb \sr~53 (
	.dataa(!virtual_state_cdr),
	.datab(!irf_reg_0_2),
	.datac(!irf_reg_1_2),
	.datad(!MonDReg_14),
	.datae(!sr_15),
	.dataf(!break_readreg_14),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~53_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~53 .extended_lut = "off";
defparam \sr~53 .lut_mask = 64'hDEFFFFFFFFFFFFFF;
defparam \sr~53 .shared_arith = "off";

cyclonev_lcell_comb \sr~54 (
	.dataa(!virtual_state_sdr),
	.datab(!altera_internal_jtag1),
	.datac(!sr_16),
	.datad(!\DRsize.010~q ),
	.datae(!\sr~53_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~54_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~54 .extended_lut = "off";
defparam \sr~54 .lut_mask = 64'h7FBFFFFF7FBFFFFF;
defparam \sr~54 .shared_arith = "off";

endmodule

module first_nios2_system_altera_std_synchronizer_2 (
	dreg_0,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_0;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module first_nios2_system_altera_std_synchronizer_3 (
	dreg_0,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_0;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module first_nios2_system_sld_virtual_jtag_basic_1 (
	virtual_state_sdr,
	virtual_state_uir1,
	virtual_state_cdr1,
	virtual_state_udr,
	state_4,
	virtual_ir_scan_reg,
	state_3,
	state_8,
	splitter_nodes_receive_1_3)/* synthesis synthesis_greybox=1 */;
output 	virtual_state_sdr;
output 	virtual_state_uir1;
output 	virtual_state_cdr1;
output 	virtual_state_udr;
input 	state_4;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_8;
input 	splitter_nodes_receive_1_3;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \virtual_state_sdr~0 (
	.dataa(!state_4),
	.datab(!virtual_ir_scan_reg),
	.datac(!splitter_nodes_receive_1_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(virtual_state_sdr),
	.sumout(),
	.cout(),
	.shareout());
defparam \virtual_state_sdr~0 .extended_lut = "off";
defparam \virtual_state_sdr~0 .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \virtual_state_sdr~0 .shared_arith = "off";

cyclonev_lcell_comb virtual_state_uir(
	.dataa(!virtual_ir_scan_reg),
	.datab(!splitter_nodes_receive_1_3),
	.datac(!state_8),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(virtual_state_uir1),
	.sumout(),
	.cout(),
	.shareout());
defparam virtual_state_uir.extended_lut = "off";
defparam virtual_state_uir.lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam virtual_state_uir.shared_arith = "off";

cyclonev_lcell_comb virtual_state_cdr(
	.dataa(!virtual_ir_scan_reg),
	.datab(!splitter_nodes_receive_1_3),
	.datac(!state_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(virtual_state_cdr1),
	.sumout(),
	.cout(),
	.shareout());
defparam virtual_state_cdr.extended_lut = "off";
defparam virtual_state_cdr.lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam virtual_state_cdr.shared_arith = "off";

cyclonev_lcell_comb \virtual_state_udr~0 (
	.dataa(!virtual_ir_scan_reg),
	.datab(!splitter_nodes_receive_1_3),
	.datac(!state_8),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(virtual_state_udr),
	.sumout(),
	.cout(),
	.shareout());
defparam \virtual_state_udr~0 .extended_lut = "off";
defparam \virtual_state_udr~0 .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \virtual_state_udr~0 .shared_arith = "off";

endmodule

module first_nios2_system_first_nios2_system_cpu_cpu_nios2_avalon_reg (
	r_sync_rst,
	oci_single_step_mode1,
	writedata_3,
	address_0,
	address_3,
	address_2,
	address_1,
	address_8,
	address_7,
	address_6,
	address_5,
	address_4,
	Equal0,
	debugaccess,
	write,
	take_action_ocireg,
	monitor_ready,
	oci_ienable_1,
	oci_ienable_16,
	writedata_1,
	writedata_16,
	oci_reg_readdata,
	oci_reg_readdata_1,
	oci_reg_readdata1,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
output 	oci_single_step_mode1;
input 	writedata_3;
input 	address_0;
input 	address_3;
input 	address_2;
input 	address_1;
input 	address_8;
input 	address_7;
input 	address_6;
input 	address_5;
input 	address_4;
output 	Equal0;
input 	debugaccess;
input 	write;
output 	take_action_ocireg;
input 	monitor_ready;
output 	oci_ienable_1;
output 	oci_ienable_16;
input 	writedata_1;
input 	writedata_16;
output 	oci_reg_readdata;
output 	oci_reg_readdata_1;
output 	oci_reg_readdata1;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \oci_single_step_mode~0_combout ;
wire \Equal0~0_combout ;
wire \oci_ienable[1]~0_combout ;
wire \Equal1~0_combout ;
wire \take_action_oci_intr_mask_reg~0_combout ;
wire \oci_ienable[16]~1_combout ;
wire \oci_ienable[0]~q ;


dffeas oci_single_step_mode(
	.clk(clk_clk),
	.d(\oci_single_step_mode~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(oci_single_step_mode1),
	.prn(vcc));
defparam oci_single_step_mode.is_wysiwyg = "true";
defparam oci_single_step_mode.power_up = "low";

cyclonev_lcell_comb \Equal0~1 (
	.dataa(!address_0),
	.datab(!address_3),
	.datac(!address_2),
	.datad(!address_1),
	.datae(!\Equal0~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal0),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~1 .extended_lut = "off";
defparam \Equal0~1 .lut_mask = 64'hFFFEFFFFFFFEFFFF;
defparam \Equal0~1 .shared_arith = "off";

cyclonev_lcell_comb \take_action_ocireg~0 (
	.dataa(!Equal0),
	.datab(!debugaccess),
	.datac(!write),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(take_action_ocireg),
	.sumout(),
	.cout(),
	.shareout());
defparam \take_action_ocireg~0 .extended_lut = "off";
defparam \take_action_ocireg~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \take_action_ocireg~0 .shared_arith = "off";

dffeas \oci_ienable[1] (
	.clk(clk_clk),
	.d(\oci_ienable[1]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_action_oci_intr_mask_reg~0_combout ),
	.q(oci_ienable_1),
	.prn(vcc));
defparam \oci_ienable[1] .is_wysiwyg = "true";
defparam \oci_ienable[1] .power_up = "low";

dffeas \oci_ienable[16] (
	.clk(clk_clk),
	.d(\oci_ienable[16]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_action_oci_intr_mask_reg~0_combout ),
	.q(oci_ienable_16),
	.prn(vcc));
defparam \oci_ienable[16] .is_wysiwyg = "true";
defparam \oci_ienable[16] .power_up = "low";

cyclonev_lcell_comb \oci_reg_readdata~0 (
	.dataa(!\Equal1~0_combout ),
	.datab(!\oci_ienable[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(oci_reg_readdata),
	.sumout(),
	.cout(),
	.shareout());
defparam \oci_reg_readdata~0 .extended_lut = "off";
defparam \oci_reg_readdata~0 .lut_mask = 64'h7777777777777777;
defparam \oci_reg_readdata~0 .shared_arith = "off";

cyclonev_lcell_comb \oci_reg_readdata[1]~1 (
	.dataa(!Equal0),
	.datab(!monitor_ready),
	.datac(!oci_ienable_1),
	.datad(!\Equal1~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(oci_reg_readdata_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \oci_reg_readdata[1]~1 .extended_lut = "off";
defparam \oci_reg_readdata[1]~1 .lut_mask = 64'hB1FFB1FFB1FFB1FF;
defparam \oci_reg_readdata[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \oci_reg_readdata~2 (
	.dataa(!oci_ienable_16),
	.datab(!\Equal1~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(oci_reg_readdata1),
	.sumout(),
	.cout(),
	.shareout());
defparam \oci_reg_readdata~2 .extended_lut = "off";
defparam \oci_reg_readdata~2 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \oci_reg_readdata~2 .shared_arith = "off";

cyclonev_lcell_comb \oci_single_step_mode~0 (
	.dataa(!oci_single_step_mode1),
	.datab(!writedata_3),
	.datac(!take_action_ocireg),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\oci_single_step_mode~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \oci_single_step_mode~0 .extended_lut = "off";
defparam \oci_single_step_mode~0 .lut_mask = 64'h5353535353535353;
defparam \oci_single_step_mode~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~0 (
	.dataa(!address_8),
	.datab(!address_7),
	.datac(!address_6),
	.datad(!address_5),
	.datae(!address_4),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~0 .extended_lut = "off";
defparam \Equal0~0 .lut_mask = 64'hFFFFFFFDFFFFFFFD;
defparam \Equal0~0 .shared_arith = "off";

cyclonev_lcell_comb \oci_ienable[1]~0 (
	.dataa(!writedata_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\oci_ienable[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \oci_ienable[1]~0 .extended_lut = "off";
defparam \oci_ienable[1]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \oci_ienable[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal1~0 (
	.dataa(!address_0),
	.datab(!address_3),
	.datac(!address_2),
	.datad(!address_1),
	.datae(!\Equal0~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal1~0 .extended_lut = "off";
defparam \Equal1~0 .lut_mask = 64'hFFFDFFFFFFFDFFFF;
defparam \Equal1~0 .shared_arith = "off";

cyclonev_lcell_comb \take_action_oci_intr_mask_reg~0 (
	.dataa(!debugaccess),
	.datab(!write),
	.datac(!\Equal1~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\take_action_oci_intr_mask_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \take_action_oci_intr_mask_reg~0 .extended_lut = "off";
defparam \take_action_oci_intr_mask_reg~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \take_action_oci_intr_mask_reg~0 .shared_arith = "off";

cyclonev_lcell_comb \oci_ienable[16]~1 (
	.dataa(!writedata_16),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\oci_ienable[16]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \oci_ienable[16]~1 .extended_lut = "off";
defparam \oci_ienable[16]~1 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \oci_ienable[16]~1 .shared_arith = "off";

dffeas \oci_ienable[0] (
	.clk(clk_clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_action_oci_intr_mask_reg~0_combout ),
	.q(\oci_ienable[0]~q ),
	.prn(vcc));
defparam \oci_ienable[0] .is_wysiwyg = "true";
defparam \oci_ienable[0] .power_up = "low";

endmodule

module first_nios2_system_first_nios2_system_cpu_cpu_nios2_oci_break (
	break_readreg_0,
	break_readreg_1,
	break_readreg_2,
	break_readreg_20,
	break_readreg_19,
	break_readreg_3,
	break_readreg_21,
	break_readreg_18,
	break_readreg_17,
	break_readreg_16,
	break_readreg_24,
	break_readreg_4,
	break_readreg_25,
	break_readreg_26,
	break_readreg_27,
	break_readreg_22,
	break_readreg_5,
	break_readreg_28,
	break_readreg_29,
	break_readreg_30,
	break_readreg_31,
	break_readreg_23,
	break_readreg_6,
	break_readreg_15,
	break_readreg_7,
	break_readreg_8,
	break_readreg_9,
	break_readreg_13,
	break_readreg_12,
	break_readreg_10,
	break_readreg_11,
	break_readreg_14,
	ir_1,
	ir_0,
	enable_action_strobe,
	jdo_21,
	jdo_20,
	jdo_0,
	jdo_36,
	jdo_37,
	jdo_3,
	jdo_19,
	jdo_18,
	jdo_17,
	jdo_25,
	jdo_1,
	jdo_4,
	jdo_26,
	jdo_27,
	jdo_28,
	jdo_2,
	jdo_5,
	jdo_29,
	jdo_30,
	jdo_31,
	jdo_23,
	jdo_22,
	jdo_6,
	jdo_24,
	jdo_16,
	jdo_7,
	jdo_8,
	jdo_9,
	jdo_10,
	jdo_14,
	jdo_13,
	jdo_11,
	jdo_12,
	jdo_15,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	break_readreg_0;
output 	break_readreg_1;
output 	break_readreg_2;
output 	break_readreg_20;
output 	break_readreg_19;
output 	break_readreg_3;
output 	break_readreg_21;
output 	break_readreg_18;
output 	break_readreg_17;
output 	break_readreg_16;
output 	break_readreg_24;
output 	break_readreg_4;
output 	break_readreg_25;
output 	break_readreg_26;
output 	break_readreg_27;
output 	break_readreg_22;
output 	break_readreg_5;
output 	break_readreg_28;
output 	break_readreg_29;
output 	break_readreg_30;
output 	break_readreg_31;
output 	break_readreg_23;
output 	break_readreg_6;
output 	break_readreg_15;
output 	break_readreg_7;
output 	break_readreg_8;
output 	break_readreg_9;
output 	break_readreg_13;
output 	break_readreg_12;
output 	break_readreg_10;
output 	break_readreg_11;
output 	break_readreg_14;
input 	ir_1;
input 	ir_0;
input 	enable_action_strobe;
input 	jdo_21;
input 	jdo_20;
input 	jdo_0;
input 	jdo_36;
input 	jdo_37;
input 	jdo_3;
input 	jdo_19;
input 	jdo_18;
input 	jdo_17;
input 	jdo_25;
input 	jdo_1;
input 	jdo_4;
input 	jdo_26;
input 	jdo_27;
input 	jdo_28;
input 	jdo_2;
input 	jdo_5;
input 	jdo_29;
input 	jdo_30;
input 	jdo_31;
input 	jdo_23;
input 	jdo_22;
input 	jdo_6;
input 	jdo_24;
input 	jdo_16;
input 	jdo_7;
input 	jdo_8;
input 	jdo_9;
input 	jdo_10;
input 	jdo_14;
input 	jdo_13;
input 	jdo_11;
input 	jdo_12;
input 	jdo_15;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \break_readreg[19]~0_combout ;
wire \break_readreg[19]~1_combout ;


dffeas \break_readreg[0] (
	.clk(clk_clk),
	.d(jdo_0),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[19]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[19]~0_combout ),
	.q(break_readreg_0),
	.prn(vcc));
defparam \break_readreg[0] .is_wysiwyg = "true";
defparam \break_readreg[0] .power_up = "low";

dffeas \break_readreg[1] (
	.clk(clk_clk),
	.d(jdo_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[19]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[19]~0_combout ),
	.q(break_readreg_1),
	.prn(vcc));
defparam \break_readreg[1] .is_wysiwyg = "true";
defparam \break_readreg[1] .power_up = "low";

dffeas \break_readreg[2] (
	.clk(clk_clk),
	.d(jdo_2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[19]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[19]~0_combout ),
	.q(break_readreg_2),
	.prn(vcc));
defparam \break_readreg[2] .is_wysiwyg = "true";
defparam \break_readreg[2] .power_up = "low";

dffeas \break_readreg[20] (
	.clk(clk_clk),
	.d(jdo_20),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[19]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[19]~0_combout ),
	.q(break_readreg_20),
	.prn(vcc));
defparam \break_readreg[20] .is_wysiwyg = "true";
defparam \break_readreg[20] .power_up = "low";

dffeas \break_readreg[19] (
	.clk(clk_clk),
	.d(jdo_19),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[19]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[19]~0_combout ),
	.q(break_readreg_19),
	.prn(vcc));
defparam \break_readreg[19] .is_wysiwyg = "true";
defparam \break_readreg[19] .power_up = "low";

dffeas \break_readreg[3] (
	.clk(clk_clk),
	.d(jdo_3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[19]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[19]~0_combout ),
	.q(break_readreg_3),
	.prn(vcc));
defparam \break_readreg[3] .is_wysiwyg = "true";
defparam \break_readreg[3] .power_up = "low";

dffeas \break_readreg[21] (
	.clk(clk_clk),
	.d(jdo_21),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[19]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[19]~0_combout ),
	.q(break_readreg_21),
	.prn(vcc));
defparam \break_readreg[21] .is_wysiwyg = "true";
defparam \break_readreg[21] .power_up = "low";

dffeas \break_readreg[18] (
	.clk(clk_clk),
	.d(jdo_18),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[19]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[19]~0_combout ),
	.q(break_readreg_18),
	.prn(vcc));
defparam \break_readreg[18] .is_wysiwyg = "true";
defparam \break_readreg[18] .power_up = "low";

dffeas \break_readreg[17] (
	.clk(clk_clk),
	.d(jdo_17),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[19]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[19]~0_combout ),
	.q(break_readreg_17),
	.prn(vcc));
defparam \break_readreg[17] .is_wysiwyg = "true";
defparam \break_readreg[17] .power_up = "low";

dffeas \break_readreg[16] (
	.clk(clk_clk),
	.d(jdo_16),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[19]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[19]~0_combout ),
	.q(break_readreg_16),
	.prn(vcc));
defparam \break_readreg[16] .is_wysiwyg = "true";
defparam \break_readreg[16] .power_up = "low";

dffeas \break_readreg[24] (
	.clk(clk_clk),
	.d(jdo_24),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[19]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[19]~0_combout ),
	.q(break_readreg_24),
	.prn(vcc));
defparam \break_readreg[24] .is_wysiwyg = "true";
defparam \break_readreg[24] .power_up = "low";

dffeas \break_readreg[4] (
	.clk(clk_clk),
	.d(jdo_4),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[19]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[19]~0_combout ),
	.q(break_readreg_4),
	.prn(vcc));
defparam \break_readreg[4] .is_wysiwyg = "true";
defparam \break_readreg[4] .power_up = "low";

dffeas \break_readreg[25] (
	.clk(clk_clk),
	.d(jdo_25),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[19]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[19]~0_combout ),
	.q(break_readreg_25),
	.prn(vcc));
defparam \break_readreg[25] .is_wysiwyg = "true";
defparam \break_readreg[25] .power_up = "low";

dffeas \break_readreg[26] (
	.clk(clk_clk),
	.d(jdo_26),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[19]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[19]~0_combout ),
	.q(break_readreg_26),
	.prn(vcc));
defparam \break_readreg[26] .is_wysiwyg = "true";
defparam \break_readreg[26] .power_up = "low";

dffeas \break_readreg[27] (
	.clk(clk_clk),
	.d(jdo_27),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[19]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[19]~0_combout ),
	.q(break_readreg_27),
	.prn(vcc));
defparam \break_readreg[27] .is_wysiwyg = "true";
defparam \break_readreg[27] .power_up = "low";

dffeas \break_readreg[22] (
	.clk(clk_clk),
	.d(jdo_22),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[19]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[19]~0_combout ),
	.q(break_readreg_22),
	.prn(vcc));
defparam \break_readreg[22] .is_wysiwyg = "true";
defparam \break_readreg[22] .power_up = "low";

dffeas \break_readreg[5] (
	.clk(clk_clk),
	.d(jdo_5),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[19]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[19]~0_combout ),
	.q(break_readreg_5),
	.prn(vcc));
defparam \break_readreg[5] .is_wysiwyg = "true";
defparam \break_readreg[5] .power_up = "low";

dffeas \break_readreg[28] (
	.clk(clk_clk),
	.d(jdo_28),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[19]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[19]~0_combout ),
	.q(break_readreg_28),
	.prn(vcc));
defparam \break_readreg[28] .is_wysiwyg = "true";
defparam \break_readreg[28] .power_up = "low";

dffeas \break_readreg[29] (
	.clk(clk_clk),
	.d(jdo_29),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[19]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[19]~0_combout ),
	.q(break_readreg_29),
	.prn(vcc));
defparam \break_readreg[29] .is_wysiwyg = "true";
defparam \break_readreg[29] .power_up = "low";

dffeas \break_readreg[30] (
	.clk(clk_clk),
	.d(jdo_30),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[19]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[19]~0_combout ),
	.q(break_readreg_30),
	.prn(vcc));
defparam \break_readreg[30] .is_wysiwyg = "true";
defparam \break_readreg[30] .power_up = "low";

dffeas \break_readreg[31] (
	.clk(clk_clk),
	.d(jdo_31),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[19]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[19]~0_combout ),
	.q(break_readreg_31),
	.prn(vcc));
defparam \break_readreg[31] .is_wysiwyg = "true";
defparam \break_readreg[31] .power_up = "low";

dffeas \break_readreg[23] (
	.clk(clk_clk),
	.d(jdo_23),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[19]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[19]~0_combout ),
	.q(break_readreg_23),
	.prn(vcc));
defparam \break_readreg[23] .is_wysiwyg = "true";
defparam \break_readreg[23] .power_up = "low";

dffeas \break_readreg[6] (
	.clk(clk_clk),
	.d(jdo_6),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[19]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[19]~0_combout ),
	.q(break_readreg_6),
	.prn(vcc));
defparam \break_readreg[6] .is_wysiwyg = "true";
defparam \break_readreg[6] .power_up = "low";

dffeas \break_readreg[15] (
	.clk(clk_clk),
	.d(jdo_15),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[19]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[19]~0_combout ),
	.q(break_readreg_15),
	.prn(vcc));
defparam \break_readreg[15] .is_wysiwyg = "true";
defparam \break_readreg[15] .power_up = "low";

dffeas \break_readreg[7] (
	.clk(clk_clk),
	.d(jdo_7),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[19]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[19]~0_combout ),
	.q(break_readreg_7),
	.prn(vcc));
defparam \break_readreg[7] .is_wysiwyg = "true";
defparam \break_readreg[7] .power_up = "low";

dffeas \break_readreg[8] (
	.clk(clk_clk),
	.d(jdo_8),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[19]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[19]~0_combout ),
	.q(break_readreg_8),
	.prn(vcc));
defparam \break_readreg[8] .is_wysiwyg = "true";
defparam \break_readreg[8] .power_up = "low";

dffeas \break_readreg[9] (
	.clk(clk_clk),
	.d(jdo_9),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[19]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[19]~0_combout ),
	.q(break_readreg_9),
	.prn(vcc));
defparam \break_readreg[9] .is_wysiwyg = "true";
defparam \break_readreg[9] .power_up = "low";

dffeas \break_readreg[13] (
	.clk(clk_clk),
	.d(jdo_13),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[19]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[19]~0_combout ),
	.q(break_readreg_13),
	.prn(vcc));
defparam \break_readreg[13] .is_wysiwyg = "true";
defparam \break_readreg[13] .power_up = "low";

dffeas \break_readreg[12] (
	.clk(clk_clk),
	.d(jdo_12),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[19]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[19]~0_combout ),
	.q(break_readreg_12),
	.prn(vcc));
defparam \break_readreg[12] .is_wysiwyg = "true";
defparam \break_readreg[12] .power_up = "low";

dffeas \break_readreg[10] (
	.clk(clk_clk),
	.d(jdo_10),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[19]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[19]~0_combout ),
	.q(break_readreg_10),
	.prn(vcc));
defparam \break_readreg[10] .is_wysiwyg = "true";
defparam \break_readreg[10] .power_up = "low";

dffeas \break_readreg[11] (
	.clk(clk_clk),
	.d(jdo_11),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[19]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[19]~0_combout ),
	.q(break_readreg_11),
	.prn(vcc));
defparam \break_readreg[11] .is_wysiwyg = "true";
defparam \break_readreg[11] .power_up = "low";

dffeas \break_readreg[14] (
	.clk(clk_clk),
	.d(jdo_14),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[19]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[19]~0_combout ),
	.q(break_readreg_14),
	.prn(vcc));
defparam \break_readreg[14] .is_wysiwyg = "true";
defparam \break_readreg[14] .power_up = "low";

cyclonev_lcell_comb \break_readreg[19]~0 (
	.dataa(!ir_1),
	.datab(!ir_0),
	.datac(!enable_action_strobe),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\break_readreg[19]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \break_readreg[19]~0 .extended_lut = "off";
defparam \break_readreg[19]~0 .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \break_readreg[19]~0 .shared_arith = "off";

cyclonev_lcell_comb \break_readreg[19]~1 (
	.dataa(!jdo_36),
	.datab(!jdo_37),
	.datac(!\break_readreg[19]~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\break_readreg[19]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \break_readreg[19]~1 .extended_lut = "off";
defparam \break_readreg[19]~1 .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \break_readreg[19]~1 .shared_arith = "off";

endmodule

module first_nios2_system_first_nios2_system_cpu_cpu_nios2_oci_debug (
	r_sync_rst,
	jtag_break1,
	take_action_ocireg,
	jdo_34,
	jdo_35,
	take_action_ocimem_a,
	take_action_ocimem_a1,
	jdo_21,
	jdo_20,
	monitor_ready1,
	jdo_19,
	jdo_18,
	jdo_25,
	writedata_0,
	writedata_1,
	monitor_error1,
	jdo_23,
	jdo_24,
	monitor_go1,
	resetlatch1,
	state_1,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
output 	jtag_break1;
input 	take_action_ocireg;
input 	jdo_34;
input 	jdo_35;
input 	take_action_ocimem_a;
input 	take_action_ocimem_a1;
input 	jdo_21;
input 	jdo_20;
output 	monitor_ready1;
input 	jdo_19;
input 	jdo_18;
input 	jdo_25;
input 	writedata_0;
input 	writedata_1;
output 	monitor_error1;
input 	jdo_23;
input 	jdo_24;
output 	monitor_go1;
output 	resetlatch1;
input 	state_1;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \the_altera_std_synchronizer|dreg[0]~q ;
wire \break_on_reset~0_combout ;
wire \break_on_reset~q ;
wire \jtag_break~0_combout ;
wire \monitor_ready~0_combout ;
wire \monitor_error~0_combout ;
wire \monitor_go~0_combout ;
wire \resetlatch~0_combout ;


first_nios2_system_altera_std_synchronizer_4 the_altera_std_synchronizer(
	.din(r_sync_rst),
	.dreg_0(\the_altera_std_synchronizer|dreg[0]~q ),
	.clk(clk_clk));

dffeas jtag_break(
	.clk(clk_clk),
	.d(\jtag_break~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(jtag_break1),
	.prn(vcc));
defparam jtag_break.is_wysiwyg = "true";
defparam jtag_break.power_up = "low";

dffeas monitor_ready(
	.clk(clk_clk),
	.d(\monitor_ready~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(monitor_ready1),
	.prn(vcc));
defparam monitor_ready.is_wysiwyg = "true";
defparam monitor_ready.power_up = "low";

dffeas monitor_error(
	.clk(clk_clk),
	.d(\monitor_error~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(monitor_error1),
	.prn(vcc));
defparam monitor_error.is_wysiwyg = "true";
defparam monitor_error.power_up = "low";

dffeas monitor_go(
	.clk(clk_clk),
	.d(\monitor_go~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(monitor_go1),
	.prn(vcc));
defparam monitor_go.is_wysiwyg = "true";
defparam monitor_go.power_up = "low";

dffeas resetlatch(
	.clk(clk_clk),
	.d(\resetlatch~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(resetlatch1),
	.prn(vcc));
defparam resetlatch.is_wysiwyg = "true";
defparam resetlatch.power_up = "low";

cyclonev_lcell_comb \break_on_reset~0 (
	.dataa(!take_action_ocimem_a1),
	.datab(!\break_on_reset~q ),
	.datac(!jdo_19),
	.datad(!jdo_18),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\break_on_reset~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \break_on_reset~0 .extended_lut = "off";
defparam \break_on_reset~0 .lut_mask = 64'hBF1FBF1FBF1FBF1F;
defparam \break_on_reset~0 .shared_arith = "off";

dffeas break_on_reset(
	.clk(clk_clk),
	.d(\break_on_reset~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\break_on_reset~q ),
	.prn(vcc));
defparam break_on_reset.is_wysiwyg = "true";
defparam break_on_reset.power_up = "low";

cyclonev_lcell_comb \jtag_break~0 (
	.dataa(!jtag_break1),
	.datab(!take_action_ocimem_a1),
	.datac(!jdo_21),
	.datad(!jdo_20),
	.datae(!\break_on_reset~q ),
	.dataf(!\the_altera_std_synchronizer|dreg[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\jtag_break~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \jtag_break~0 .extended_lut = "off";
defparam \jtag_break~0 .lut_mask = 64'hFF7FFFFFFFDFFFFF;
defparam \jtag_break~0 .shared_arith = "off";

cyclonev_lcell_comb \monitor_ready~0 (
	.dataa(!take_action_ocireg),
	.datab(!take_action_ocimem_a1),
	.datac(!monitor_ready1),
	.datad(!jdo_25),
	.datae(!writedata_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\monitor_ready~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \monitor_ready~0 .extended_lut = "off";
defparam \monitor_ready~0 .lut_mask = 64'hFFDFFFFFFFDFFFFF;
defparam \monitor_ready~0 .shared_arith = "off";

cyclonev_lcell_comb \monitor_error~0 (
	.dataa(!take_action_ocireg),
	.datab(!take_action_ocimem_a1),
	.datac(!jdo_25),
	.datad(!writedata_1),
	.datae(!monitor_error1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\monitor_error~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \monitor_error~0 .extended_lut = "off";
defparam \monitor_error~0 .lut_mask = 64'hFDFFFFFFFDFFFFFF;
defparam \monitor_error~0 .shared_arith = "off";

cyclonev_lcell_comb \monitor_go~0 (
	.dataa(!jdo_34),
	.datab(!jdo_35),
	.datac(!take_action_ocimem_a),
	.datad(!jdo_23),
	.datae(!monitor_go1),
	.dataf(!state_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\monitor_go~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \monitor_go~0 .extended_lut = "off";
defparam \monitor_go~0 .lut_mask = 64'hFFFFFFFFDFFFFFFF;
defparam \monitor_go~0 .shared_arith = "off";

cyclonev_lcell_comb \resetlatch~0 (
	.dataa(!take_action_ocimem_a1),
	.datab(!\the_altera_std_synchronizer|dreg[0]~q ),
	.datac(!jdo_24),
	.datad(!resetlatch1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\resetlatch~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \resetlatch~0 .extended_lut = "off";
defparam \resetlatch~0 .lut_mask = 64'hFBFFFBFFFBFFFBFF;
defparam \resetlatch~0 .shared_arith = "off";

endmodule

module first_nios2_system_altera_std_synchronizer_4 (
	din,
	dreg_0,
	clk)/* synthesis synthesis_greybox=1 */;
input 	din;
output 	dreg_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module first_nios2_system_first_nios2_system_cpu_cpu_nios2_ocimem (
	q_a_0,
	MonDReg_2,
	q_a_1,
	MonDReg_20,
	MonDReg_19,
	q_a_2,
	MonDReg_21,
	q_a_20,
	q_a_19,
	MonDReg_17,
	MonDReg_16,
	MonDReg_24,
	q_a_3,
	MonDReg_25,
	MonDReg_26,
	MonDReg_27,
	q_a_21,
	q_a_18,
	q_a_17,
	q_a_16,
	q_a_4,
	q_a_5,
	q_a_6,
	q_a_7,
	q_a_24,
	q_a_25,
	q_a_26,
	MonDReg_28,
	q_a_27,
	MonDReg_30,
	MonDReg_31,
	q_a_22,
	q_a_23,
	q_a_31,
	q_a_11,
	q_a_28,
	q_a_10,
	q_a_8,
	q_a_9,
	q_a_30,
	q_a_15,
	q_a_12,
	q_a_13,
	q_a_14,
	q_a_29,
	MonDReg_23,
	MonDReg_6,
	MonDReg_7,
	MonDReg_11,
	MonDReg_10,
	MonDReg_9,
	MonDReg_13,
	MonDReg_14,
	waitrequest1,
	MonDReg_0,
	writedata_3,
	address_0,
	address_3,
	address_2,
	address_1,
	address_8,
	address_7,
	address_6,
	address_5,
	address_4,
	debugaccess,
	write,
	jdo_34,
	jdo_35,
	take_action_ocimem_a,
	take_no_action_ocimem_a,
	take_action_ocimem_a1,
	jdo_21,
	jdo_20,
	read,
	MonDReg_1,
	jdo_3,
	jdo_19,
	jdo_18,
	jdo_17,
	jdo_25,
	writedata_0,
	jdo_4,
	jdo_26,
	jdo_27,
	jdo_28,
	r_early_rst,
	byteenable_0,
	writedata_1,
	writedata_16,
	MonDReg_3,
	jdo_5,
	jdo_29,
	jdo_30,
	jdo_31,
	jdo_32,
	jdo_33,
	jdo_23,
	jdo_22,
	MonDReg_18,
	MonDReg_4,
	jdo_6,
	writedata_2,
	MonDReg_22,
	jdo_24,
	writedata_20,
	byteenable_2,
	writedata_19,
	jdo_16,
	MonDReg_5,
	jdo_7,
	MonDReg_29,
	writedata_21,
	writedata_18,
	writedata_17,
	writedata_4,
	writedata_5,
	writedata_6,
	writedata_7,
	writedata_24,
	byteenable_3,
	jdo_8,
	writedata_25,
	writedata_26,
	writedata_27,
	writedata_22,
	writedata_23,
	writedata_31,
	writedata_11,
	byteenable_1,
	writedata_28,
	writedata_10,
	MonDReg_8,
	writedata_8,
	writedata_9,
	writedata_30,
	MonDReg_15,
	writedata_15,
	MonDReg_12,
	writedata_12,
	writedata_13,
	writedata_14,
	writedata_29,
	jdo_9,
	jdo_10,
	jdo_14,
	jdo_13,
	jdo_11,
	jdo_12,
	jdo_15,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	q_a_0;
output 	MonDReg_2;
output 	q_a_1;
output 	MonDReg_20;
output 	MonDReg_19;
output 	q_a_2;
output 	MonDReg_21;
output 	q_a_20;
output 	q_a_19;
output 	MonDReg_17;
output 	MonDReg_16;
output 	MonDReg_24;
output 	q_a_3;
output 	MonDReg_25;
output 	MonDReg_26;
output 	MonDReg_27;
output 	q_a_21;
output 	q_a_18;
output 	q_a_17;
output 	q_a_16;
output 	q_a_4;
output 	q_a_5;
output 	q_a_6;
output 	q_a_7;
output 	q_a_24;
output 	q_a_25;
output 	q_a_26;
output 	MonDReg_28;
output 	q_a_27;
output 	MonDReg_30;
output 	MonDReg_31;
output 	q_a_22;
output 	q_a_23;
output 	q_a_31;
output 	q_a_11;
output 	q_a_28;
output 	q_a_10;
output 	q_a_8;
output 	q_a_9;
output 	q_a_30;
output 	q_a_15;
output 	q_a_12;
output 	q_a_13;
output 	q_a_14;
output 	q_a_29;
output 	MonDReg_23;
output 	MonDReg_6;
output 	MonDReg_7;
output 	MonDReg_11;
output 	MonDReg_10;
output 	MonDReg_9;
output 	MonDReg_13;
output 	MonDReg_14;
output 	waitrequest1;
output 	MonDReg_0;
input 	writedata_3;
input 	address_0;
input 	address_3;
input 	address_2;
input 	address_1;
input 	address_8;
input 	address_7;
input 	address_6;
input 	address_5;
input 	address_4;
input 	debugaccess;
input 	write;
input 	jdo_34;
input 	jdo_35;
input 	take_action_ocimem_a;
input 	take_no_action_ocimem_a;
input 	take_action_ocimem_a1;
input 	jdo_21;
input 	jdo_20;
input 	read;
output 	MonDReg_1;
input 	jdo_3;
input 	jdo_19;
input 	jdo_18;
input 	jdo_17;
input 	jdo_25;
input 	writedata_0;
input 	jdo_4;
input 	jdo_26;
input 	jdo_27;
input 	jdo_28;
input 	r_early_rst;
input 	byteenable_0;
input 	writedata_1;
input 	writedata_16;
output 	MonDReg_3;
input 	jdo_5;
input 	jdo_29;
input 	jdo_30;
input 	jdo_31;
input 	jdo_32;
input 	jdo_33;
input 	jdo_23;
input 	jdo_22;
output 	MonDReg_18;
output 	MonDReg_4;
input 	jdo_6;
input 	writedata_2;
output 	MonDReg_22;
input 	jdo_24;
input 	writedata_20;
input 	byteenable_2;
input 	writedata_19;
input 	jdo_16;
output 	MonDReg_5;
input 	jdo_7;
output 	MonDReg_29;
input 	writedata_21;
input 	writedata_18;
input 	writedata_17;
input 	writedata_4;
input 	writedata_5;
input 	writedata_6;
input 	writedata_7;
input 	writedata_24;
input 	byteenable_3;
input 	jdo_8;
input 	writedata_25;
input 	writedata_26;
input 	writedata_27;
input 	writedata_22;
input 	writedata_23;
input 	writedata_31;
input 	writedata_11;
input 	byteenable_1;
input 	writedata_28;
input 	writedata_10;
output 	MonDReg_8;
input 	writedata_8;
input 	writedata_9;
input 	writedata_30;
output 	MonDReg_15;
input 	writedata_15;
output 	MonDReg_12;
input 	writedata_12;
input 	writedata_13;
input 	writedata_14;
input 	writedata_29;
input 	jdo_9;
input 	jdo_10;
input 	jdo_14;
input 	jdo_13;
input 	jdo_11;
input 	jdo_12;
input 	jdo_15;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \jtag_ram_wr~q ;
wire \ociram_wr_en~0_combout ;
wire \ociram_reset_req~combout ;
wire \ociram_wr_data[0]~0_combout ;
wire \ociram_addr[0]~0_combout ;
wire \ociram_addr[1]~1_combout ;
wire \ociram_addr[2]~2_combout ;
wire \ociram_addr[3]~3_combout ;
wire \ociram_addr[4]~4_combout ;
wire \ociram_addr[5]~5_combout ;
wire \ociram_addr[6]~6_combout ;
wire \ociram_addr[7]~7_combout ;
wire \ociram_byteenable[0]~0_combout ;
wire \ociram_wr_data[1]~1_combout ;
wire \jtag_ram_wr~0_combout ;
wire \ociram_wr_data[2]~2_combout ;
wire \ociram_wr_data[20]~3_combout ;
wire \ociram_byteenable[2]~1_combout ;
wire \ociram_wr_data[19]~4_combout ;
wire \ociram_wr_data[3]~5_combout ;
wire \ociram_wr_data[21]~6_combout ;
wire \ociram_wr_data[18]~7_combout ;
wire \ociram_wr_data[17]~8_combout ;
wire \ociram_wr_data[16]~9_combout ;
wire \ociram_wr_data[4]~10_combout ;
wire \ociram_wr_data[5]~11_combout ;
wire \ociram_wr_data[6]~12_combout ;
wire \ociram_wr_data[7]~13_combout ;
wire \ociram_wr_data[24]~14_combout ;
wire \ociram_byteenable[3]~2_combout ;
wire \ociram_wr_data[25]~15_combout ;
wire \ociram_wr_data[26]~16_combout ;
wire \ociram_wr_data[27]~17_combout ;
wire \ociram_wr_data[22]~18_combout ;
wire \ociram_wr_data[23]~19_combout ;
wire \ociram_wr_data[31]~20_combout ;
wire \ociram_wr_data[11]~21_combout ;
wire \ociram_byteenable[1]~3_combout ;
wire \ociram_wr_data[28]~22_combout ;
wire \ociram_wr_data[10]~23_combout ;
wire \ociram_wr_data[8]~24_combout ;
wire \ociram_wr_data[9]~25_combout ;
wire \ociram_wr_data[30]~26_combout ;
wire \ociram_wr_data[15]~27_combout ;
wire \ociram_wr_data[12]~28_combout ;
wire \ociram_wr_data[13]~29_combout ;
wire \ociram_wr_data[14]~30_combout ;
wire \ociram_wr_data[29]~31_combout ;
wire \Add0~1_wirecell_combout ;
wire \MonAReg[10]~q ;
wire \Add0~5_sumout ;
wire \MonAReg[2]~q ;
wire \Add0~6 ;
wire \Add0~9_sumout ;
wire \MonAReg[3]~q ;
wire \Add0~10 ;
wire \Add0~13_sumout ;
wire \MonAReg[4]~q ;
wire \Add0~14 ;
wire \Add0~21_sumout ;
wire \MonAReg[5]~q ;
wire \Add0~22 ;
wire \Add0~25_sumout ;
wire \MonAReg[6]~q ;
wire \Add0~26 ;
wire \Add0~29_sumout ;
wire \MonAReg[7]~q ;
wire \Add0~30 ;
wire \Add0~33_sumout ;
wire \MonAReg[8]~q ;
wire \Add0~34 ;
wire \Add0~17_sumout ;
wire \MonAReg[9]~q ;
wire \Add0~18 ;
wire \Add0~1_sumout ;
wire \jtag_ram_rd~0_combout ;
wire \MonDReg[8]~0_combout ;
wire \jtag_ram_rd~q ;
wire \jtag_ram_rd_d1~q ;
wire \MonDReg[8]~1_combout ;
wire \jtag_rd~q ;
wire \jtag_rd_d1~q ;
wire \MonDReg[0]~2_combout ;
wire \jtag_ram_access~0_combout ;
wire \jtag_ram_access~q ;
wire \waitrequest~0_combout ;
wire \avalon_ociram_readdata_ready~0_combout ;
wire \avalon_ociram_readdata_ready~q ;
wire \waitrequest~1_combout ;
wire \MonDReg~16_combout ;
wire \Equal0~0_combout ;
wire \MonDReg~3_combout ;
wire \MonDReg~4_combout ;
wire \MonDReg~5_combout ;
wire \MonDReg~6_combout ;
wire \MonDReg~7_combout ;
wire \MonDReg~8_combout ;
wire \MonDReg~9_combout ;
wire \Equal0~1_combout ;
wire \MonDReg~10_combout ;
wire \MonDReg~11_combout ;
wire \MonDReg~15_combout ;
wire \MonDReg~14_combout ;
wire \MonDReg~12_combout ;
wire \MonDReg~13_combout ;


first_nios2_system_first_nios2_system_cpu_cpu_ociram_sp_ram_module first_nios2_system_cpu_cpu_ociram_sp_ram(
	.q_a_0(q_a_0),
	.q_a_1(q_a_1),
	.q_a_2(q_a_2),
	.q_a_20(q_a_20),
	.q_a_19(q_a_19),
	.q_a_3(q_a_3),
	.q_a_21(q_a_21),
	.q_a_18(q_a_18),
	.q_a_17(q_a_17),
	.q_a_16(q_a_16),
	.q_a_4(q_a_4),
	.q_a_5(q_a_5),
	.q_a_6(q_a_6),
	.q_a_7(q_a_7),
	.q_a_24(q_a_24),
	.q_a_25(q_a_25),
	.q_a_26(q_a_26),
	.q_a_27(q_a_27),
	.q_a_22(q_a_22),
	.q_a_23(q_a_23),
	.q_a_31(q_a_31),
	.q_a_11(q_a_11),
	.q_a_28(q_a_28),
	.q_a_10(q_a_10),
	.q_a_8(q_a_8),
	.q_a_9(q_a_9),
	.q_a_30(q_a_30),
	.q_a_15(q_a_15),
	.q_a_12(q_a_12),
	.q_a_13(q_a_13),
	.q_a_14(q_a_14),
	.q_a_29(q_a_29),
	.ociram_wr_en(\ociram_wr_en~0_combout ),
	.ociram_reset_req(\ociram_reset_req~combout ),
	.ociram_wr_data_0(\ociram_wr_data[0]~0_combout ),
	.ociram_addr_0(\ociram_addr[0]~0_combout ),
	.ociram_addr_1(\ociram_addr[1]~1_combout ),
	.ociram_addr_2(\ociram_addr[2]~2_combout ),
	.ociram_addr_3(\ociram_addr[3]~3_combout ),
	.ociram_addr_4(\ociram_addr[4]~4_combout ),
	.ociram_addr_5(\ociram_addr[5]~5_combout ),
	.ociram_addr_6(\ociram_addr[6]~6_combout ),
	.ociram_addr_7(\ociram_addr[7]~7_combout ),
	.ociram_byteenable_0(\ociram_byteenable[0]~0_combout ),
	.ociram_wr_data_1(\ociram_wr_data[1]~1_combout ),
	.ociram_wr_data_2(\ociram_wr_data[2]~2_combout ),
	.ociram_wr_data_20(\ociram_wr_data[20]~3_combout ),
	.ociram_byteenable_2(\ociram_byteenable[2]~1_combout ),
	.ociram_wr_data_19(\ociram_wr_data[19]~4_combout ),
	.ociram_wr_data_3(\ociram_wr_data[3]~5_combout ),
	.ociram_wr_data_21(\ociram_wr_data[21]~6_combout ),
	.ociram_wr_data_18(\ociram_wr_data[18]~7_combout ),
	.ociram_wr_data_17(\ociram_wr_data[17]~8_combout ),
	.ociram_wr_data_16(\ociram_wr_data[16]~9_combout ),
	.ociram_wr_data_4(\ociram_wr_data[4]~10_combout ),
	.ociram_wr_data_5(\ociram_wr_data[5]~11_combout ),
	.ociram_wr_data_6(\ociram_wr_data[6]~12_combout ),
	.ociram_wr_data_7(\ociram_wr_data[7]~13_combout ),
	.ociram_wr_data_24(\ociram_wr_data[24]~14_combout ),
	.ociram_byteenable_3(\ociram_byteenable[3]~2_combout ),
	.ociram_wr_data_25(\ociram_wr_data[25]~15_combout ),
	.ociram_wr_data_26(\ociram_wr_data[26]~16_combout ),
	.ociram_wr_data_27(\ociram_wr_data[27]~17_combout ),
	.ociram_wr_data_22(\ociram_wr_data[22]~18_combout ),
	.ociram_wr_data_23(\ociram_wr_data[23]~19_combout ),
	.ociram_wr_data_31(\ociram_wr_data[31]~20_combout ),
	.ociram_wr_data_11(\ociram_wr_data[11]~21_combout ),
	.ociram_byteenable_1(\ociram_byteenable[1]~3_combout ),
	.ociram_wr_data_28(\ociram_wr_data[28]~22_combout ),
	.ociram_wr_data_10(\ociram_wr_data[10]~23_combout ),
	.ociram_wr_data_8(\ociram_wr_data[8]~24_combout ),
	.ociram_wr_data_9(\ociram_wr_data[9]~25_combout ),
	.ociram_wr_data_30(\ociram_wr_data[30]~26_combout ),
	.ociram_wr_data_15(\ociram_wr_data[15]~27_combout ),
	.ociram_wr_data_12(\ociram_wr_data[12]~28_combout ),
	.ociram_wr_data_13(\ociram_wr_data[13]~29_combout ),
	.ociram_wr_data_14(\ociram_wr_data[14]~30_combout ),
	.ociram_wr_data_29(\ociram_wr_data[29]~31_combout ),
	.clk_clk(clk_clk));

dffeas jtag_ram_wr(
	.clk(clk_clk),
	.d(\jtag_ram_wr~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!take_no_action_ocimem_a),
	.q(\jtag_ram_wr~q ),
	.prn(vcc));
defparam jtag_ram_wr.is_wysiwyg = "true";
defparam jtag_ram_wr.power_up = "low";

cyclonev_lcell_comb \ociram_wr_en~0 (
	.dataa(!address_8),
	.datab(!debugaccess),
	.datac(!write),
	.datad(!\jtag_ram_access~q ),
	.datae(!\jtag_ram_wr~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_en~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_en~0 .extended_lut = "off";
defparam \ociram_wr_en~0 .lut_mask = 64'hAF3FFFFFAF3FFFFF;
defparam \ociram_wr_en~0 .shared_arith = "off";

cyclonev_lcell_comb ociram_reset_req(
	.dataa(!\jtag_ram_access~q ),
	.datab(!r_early_rst),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_reset_req~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam ociram_reset_req.extended_lut = "off";
defparam ociram_reset_req.lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam ociram_reset_req.shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[0]~0 (
	.dataa(!MonDReg_0),
	.datab(!\jtag_ram_access~q ),
	.datac(!writedata_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[0]~0 .extended_lut = "off";
defparam \ociram_wr_data[0]~0 .lut_mask = 64'h4747474747474747;
defparam \ociram_wr_data[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \ociram_addr[0]~0 (
	.dataa(!address_0),
	.datab(!\jtag_ram_access~q ),
	.datac(!\MonAReg[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_addr[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_addr[0]~0 .extended_lut = "off";
defparam \ociram_addr[0]~0 .lut_mask = 64'h4747474747474747;
defparam \ociram_addr[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \ociram_addr[1]~1 (
	.dataa(!address_1),
	.datab(!\jtag_ram_access~q ),
	.datac(!\MonAReg[3]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_addr[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_addr[1]~1 .extended_lut = "off";
defparam \ociram_addr[1]~1 .lut_mask = 64'h4747474747474747;
defparam \ociram_addr[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \ociram_addr[2]~2 (
	.dataa(!address_2),
	.datab(!\jtag_ram_access~q ),
	.datac(!\MonAReg[4]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_addr[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_addr[2]~2 .extended_lut = "off";
defparam \ociram_addr[2]~2 .lut_mask = 64'h4747474747474747;
defparam \ociram_addr[2]~2 .shared_arith = "off";

cyclonev_lcell_comb \ociram_addr[3]~3 (
	.dataa(!address_3),
	.datab(!\jtag_ram_access~q ),
	.datac(!\MonAReg[5]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_addr[3]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_addr[3]~3 .extended_lut = "off";
defparam \ociram_addr[3]~3 .lut_mask = 64'h4747474747474747;
defparam \ociram_addr[3]~3 .shared_arith = "off";

cyclonev_lcell_comb \ociram_addr[4]~4 (
	.dataa(!address_4),
	.datab(!\jtag_ram_access~q ),
	.datac(!\MonAReg[6]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_addr[4]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_addr[4]~4 .extended_lut = "off";
defparam \ociram_addr[4]~4 .lut_mask = 64'h4747474747474747;
defparam \ociram_addr[4]~4 .shared_arith = "off";

cyclonev_lcell_comb \ociram_addr[5]~5 (
	.dataa(!address_5),
	.datab(!\jtag_ram_access~q ),
	.datac(!\MonAReg[7]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_addr[5]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_addr[5]~5 .extended_lut = "off";
defparam \ociram_addr[5]~5 .lut_mask = 64'h4747474747474747;
defparam \ociram_addr[5]~5 .shared_arith = "off";

cyclonev_lcell_comb \ociram_addr[6]~6 (
	.dataa(!address_6),
	.datab(!\jtag_ram_access~q ),
	.datac(!\MonAReg[8]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_addr[6]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_addr[6]~6 .extended_lut = "off";
defparam \ociram_addr[6]~6 .lut_mask = 64'h4747474747474747;
defparam \ociram_addr[6]~6 .shared_arith = "off";

cyclonev_lcell_comb \ociram_addr[7]~7 (
	.dataa(!address_7),
	.datab(!\jtag_ram_access~q ),
	.datac(!\MonAReg[9]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_addr[7]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_addr[7]~7 .extended_lut = "off";
defparam \ociram_addr[7]~7 .lut_mask = 64'h4747474747474747;
defparam \ociram_addr[7]~7 .shared_arith = "off";

cyclonev_lcell_comb \ociram_byteenable[0]~0 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!byteenable_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_byteenable[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_byteenable[0]~0 .extended_lut = "off";
defparam \ociram_byteenable[0]~0 .lut_mask = 64'h7777777777777777;
defparam \ociram_byteenable[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[1]~1 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_1),
	.datac(!writedata_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[1]~1 .extended_lut = "off";
defparam \ociram_wr_data[1]~1 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \jtag_ram_wr~0 (
	.dataa(!\MonDReg[8]~0_combout ),
	.datab(!\Add0~1_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\jtag_ram_wr~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \jtag_ram_wr~0 .extended_lut = "off";
defparam \jtag_ram_wr~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \jtag_ram_wr~0 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[2]~2 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_2),
	.datac(!writedata_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[2]~2 .extended_lut = "off";
defparam \ociram_wr_data[2]~2 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[2]~2 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[20]~3 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_20),
	.datac(!writedata_20),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[20]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[20]~3 .extended_lut = "off";
defparam \ociram_wr_data[20]~3 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[20]~3 .shared_arith = "off";

cyclonev_lcell_comb \ociram_byteenable[2]~1 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!byteenable_2),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_byteenable[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_byteenable[2]~1 .extended_lut = "off";
defparam \ociram_byteenable[2]~1 .lut_mask = 64'h7777777777777777;
defparam \ociram_byteenable[2]~1 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[19]~4 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_19),
	.datac(!writedata_19),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[19]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[19]~4 .extended_lut = "off";
defparam \ociram_wr_data[19]~4 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[19]~4 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[3]~5 (
	.dataa(!writedata_3),
	.datab(!\jtag_ram_access~q ),
	.datac(!MonDReg_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[3]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[3]~5 .extended_lut = "off";
defparam \ociram_wr_data[3]~5 .lut_mask = 64'h4747474747474747;
defparam \ociram_wr_data[3]~5 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[21]~6 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_21),
	.datac(!writedata_21),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[21]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[21]~6 .extended_lut = "off";
defparam \ociram_wr_data[21]~6 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[21]~6 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[18]~7 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_18),
	.datac(!writedata_18),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[18]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[18]~7 .extended_lut = "off";
defparam \ociram_wr_data[18]~7 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[18]~7 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[17]~8 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_17),
	.datac(!writedata_17),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[17]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[17]~8 .extended_lut = "off";
defparam \ociram_wr_data[17]~8 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[17]~8 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[16]~9 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!writedata_16),
	.datac(!MonDReg_16),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[16]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[16]~9 .extended_lut = "off";
defparam \ociram_wr_data[16]~9 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[16]~9 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[4]~10 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_4),
	.datac(!writedata_4),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[4]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[4]~10 .extended_lut = "off";
defparam \ociram_wr_data[4]~10 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[4]~10 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[5]~11 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_5),
	.datac(!writedata_5),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[5]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[5]~11 .extended_lut = "off";
defparam \ociram_wr_data[5]~11 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[5]~11 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[6]~12 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_6),
	.datac(!writedata_6),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[6]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[6]~12 .extended_lut = "off";
defparam \ociram_wr_data[6]~12 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[6]~12 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[7]~13 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_7),
	.datac(!writedata_7),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[7]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[7]~13 .extended_lut = "off";
defparam \ociram_wr_data[7]~13 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[7]~13 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[24]~14 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_24),
	.datac(!writedata_24),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[24]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[24]~14 .extended_lut = "off";
defparam \ociram_wr_data[24]~14 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[24]~14 .shared_arith = "off";

cyclonev_lcell_comb \ociram_byteenable[3]~2 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!byteenable_3),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_byteenable[3]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_byteenable[3]~2 .extended_lut = "off";
defparam \ociram_byteenable[3]~2 .lut_mask = 64'h7777777777777777;
defparam \ociram_byteenable[3]~2 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[25]~15 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_25),
	.datac(!writedata_25),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[25]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[25]~15 .extended_lut = "off";
defparam \ociram_wr_data[25]~15 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[25]~15 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[26]~16 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_26),
	.datac(!writedata_26),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[26]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[26]~16 .extended_lut = "off";
defparam \ociram_wr_data[26]~16 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[26]~16 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[27]~17 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_27),
	.datac(!writedata_27),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[27]~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[27]~17 .extended_lut = "off";
defparam \ociram_wr_data[27]~17 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[27]~17 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[22]~18 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_22),
	.datac(!writedata_22),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[22]~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[22]~18 .extended_lut = "off";
defparam \ociram_wr_data[22]~18 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[22]~18 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[23]~19 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_23),
	.datac(!writedata_23),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[23]~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[23]~19 .extended_lut = "off";
defparam \ociram_wr_data[23]~19 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[23]~19 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[31]~20 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_31),
	.datac(!writedata_31),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[31]~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[31]~20 .extended_lut = "off";
defparam \ociram_wr_data[31]~20 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[31]~20 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[11]~21 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_11),
	.datac(!writedata_11),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[11]~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[11]~21 .extended_lut = "off";
defparam \ociram_wr_data[11]~21 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[11]~21 .shared_arith = "off";

cyclonev_lcell_comb \ociram_byteenable[1]~3 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!byteenable_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_byteenable[1]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_byteenable[1]~3 .extended_lut = "off";
defparam \ociram_byteenable[1]~3 .lut_mask = 64'h7777777777777777;
defparam \ociram_byteenable[1]~3 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[28]~22 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_28),
	.datac(!writedata_28),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[28]~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[28]~22 .extended_lut = "off";
defparam \ociram_wr_data[28]~22 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[28]~22 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[10]~23 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_10),
	.datac(!writedata_10),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[10]~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[10]~23 .extended_lut = "off";
defparam \ociram_wr_data[10]~23 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[10]~23 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[8]~24 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_8),
	.datac(!writedata_8),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[8]~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[8]~24 .extended_lut = "off";
defparam \ociram_wr_data[8]~24 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[8]~24 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[9]~25 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_9),
	.datac(!writedata_9),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[9]~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[9]~25 .extended_lut = "off";
defparam \ociram_wr_data[9]~25 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[9]~25 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[30]~26 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_30),
	.datac(!writedata_30),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[30]~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[30]~26 .extended_lut = "off";
defparam \ociram_wr_data[30]~26 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[30]~26 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[15]~27 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_15),
	.datac(!writedata_15),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[15]~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[15]~27 .extended_lut = "off";
defparam \ociram_wr_data[15]~27 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[15]~27 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[12]~28 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_12),
	.datac(!writedata_12),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[12]~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[12]~28 .extended_lut = "off";
defparam \ociram_wr_data[12]~28 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[12]~28 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[13]~29 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_13),
	.datac(!writedata_13),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[13]~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[13]~29 .extended_lut = "off";
defparam \ociram_wr_data[13]~29 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[13]~29 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[14]~30 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_14),
	.datac(!writedata_14),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[14]~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[14]~30 .extended_lut = "off";
defparam \ociram_wr_data[14]~30 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[14]~30 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[29]~31 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_29),
	.datac(!writedata_29),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[29]~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[29]~31 .extended_lut = "off";
defparam \ociram_wr_data[29]~31 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[29]~31 .shared_arith = "off";

dffeas \MonDReg[2] (
	.clk(clk_clk),
	.d(jdo_5),
	.asdata(q_a_2),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[8]~1_combout ),
	.sload(\MonDReg[8]~0_combout ),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_2),
	.prn(vcc));
defparam \MonDReg[2] .is_wysiwyg = "true";
defparam \MonDReg[2] .power_up = "low";

dffeas \MonDReg[20] (
	.clk(clk_clk),
	.d(jdo_23),
	.asdata(q_a_20),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[8]~1_combout ),
	.sload(\MonDReg[8]~0_combout ),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_20),
	.prn(vcc));
defparam \MonDReg[20] .is_wysiwyg = "true";
defparam \MonDReg[20] .power_up = "low";

dffeas \MonDReg[19] (
	.clk(clk_clk),
	.d(jdo_22),
	.asdata(q_a_19),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[8]~1_combout ),
	.sload(\MonDReg[8]~0_combout ),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_19),
	.prn(vcc));
defparam \MonDReg[19] .is_wysiwyg = "true";
defparam \MonDReg[19] .power_up = "low";

dffeas \MonDReg[21] (
	.clk(clk_clk),
	.d(jdo_24),
	.asdata(q_a_21),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[8]~1_combout ),
	.sload(\MonDReg[8]~0_combout ),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_21),
	.prn(vcc));
defparam \MonDReg[21] .is_wysiwyg = "true";
defparam \MonDReg[21] .power_up = "low";

dffeas \MonDReg[17] (
	.clk(clk_clk),
	.d(jdo_20),
	.asdata(q_a_17),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[8]~1_combout ),
	.sload(\MonDReg[8]~0_combout ),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_17),
	.prn(vcc));
defparam \MonDReg[17] .is_wysiwyg = "true";
defparam \MonDReg[17] .power_up = "low";

dffeas \MonDReg[16] (
	.clk(clk_clk),
	.d(jdo_19),
	.asdata(q_a_16),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[8]~1_combout ),
	.sload(\MonDReg[8]~0_combout ),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_16),
	.prn(vcc));
defparam \MonDReg[16] .is_wysiwyg = "true";
defparam \MonDReg[16] .power_up = "low";

dffeas \MonDReg[24] (
	.clk(clk_clk),
	.d(jdo_27),
	.asdata(q_a_24),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[8]~1_combout ),
	.sload(\MonDReg[8]~0_combout ),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_24),
	.prn(vcc));
defparam \MonDReg[24] .is_wysiwyg = "true";
defparam \MonDReg[24] .power_up = "low";

dffeas \MonDReg[25] (
	.clk(clk_clk),
	.d(jdo_28),
	.asdata(q_a_25),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[8]~1_combout ),
	.sload(\MonDReg[8]~0_combout ),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_25),
	.prn(vcc));
defparam \MonDReg[25] .is_wysiwyg = "true";
defparam \MonDReg[25] .power_up = "low";

dffeas \MonDReg[26] (
	.clk(clk_clk),
	.d(jdo_29),
	.asdata(q_a_26),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[8]~1_combout ),
	.sload(\MonDReg[8]~0_combout ),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_26),
	.prn(vcc));
defparam \MonDReg[26] .is_wysiwyg = "true";
defparam \MonDReg[26] .power_up = "low";

dffeas \MonDReg[27] (
	.clk(clk_clk),
	.d(jdo_30),
	.asdata(q_a_27),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[8]~1_combout ),
	.sload(\MonDReg[8]~0_combout ),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_27),
	.prn(vcc));
defparam \MonDReg[27] .is_wysiwyg = "true";
defparam \MonDReg[27] .power_up = "low";

dffeas \MonDReg[28] (
	.clk(clk_clk),
	.d(jdo_31),
	.asdata(q_a_28),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[8]~1_combout ),
	.sload(\MonDReg[8]~0_combout ),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_28),
	.prn(vcc));
defparam \MonDReg[28] .is_wysiwyg = "true";
defparam \MonDReg[28] .power_up = "low";

dffeas \MonDReg[30] (
	.clk(clk_clk),
	.d(jdo_33),
	.asdata(q_a_30),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[8]~1_combout ),
	.sload(\MonDReg[8]~0_combout ),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_30),
	.prn(vcc));
defparam \MonDReg[30] .is_wysiwyg = "true";
defparam \MonDReg[30] .power_up = "low";

dffeas \MonDReg[31] (
	.clk(clk_clk),
	.d(jdo_34),
	.asdata(q_a_31),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[8]~1_combout ),
	.sload(\MonDReg[8]~0_combout ),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_31),
	.prn(vcc));
defparam \MonDReg[31] .is_wysiwyg = "true";
defparam \MonDReg[31] .power_up = "low";

dffeas \MonDReg[23] (
	.clk(clk_clk),
	.d(jdo_26),
	.asdata(q_a_23),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[8]~1_combout ),
	.sload(\MonDReg[8]~0_combout ),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_23),
	.prn(vcc));
defparam \MonDReg[23] .is_wysiwyg = "true";
defparam \MonDReg[23] .power_up = "low";

dffeas \MonDReg[6] (
	.clk(clk_clk),
	.d(jdo_9),
	.asdata(q_a_6),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[8]~1_combout ),
	.sload(\MonDReg[8]~0_combout ),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_6),
	.prn(vcc));
defparam \MonDReg[6] .is_wysiwyg = "true";
defparam \MonDReg[6] .power_up = "low";

dffeas \MonDReg[7] (
	.clk(clk_clk),
	.d(jdo_10),
	.asdata(q_a_7),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[8]~1_combout ),
	.sload(\MonDReg[8]~0_combout ),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_7),
	.prn(vcc));
defparam \MonDReg[7] .is_wysiwyg = "true";
defparam \MonDReg[7] .power_up = "low";

dffeas \MonDReg[11] (
	.clk(clk_clk),
	.d(jdo_14),
	.asdata(q_a_11),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[8]~1_combout ),
	.sload(\MonDReg[8]~0_combout ),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_11),
	.prn(vcc));
defparam \MonDReg[11] .is_wysiwyg = "true";
defparam \MonDReg[11] .power_up = "low";

dffeas \MonDReg[10] (
	.clk(clk_clk),
	.d(jdo_13),
	.asdata(q_a_10),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[8]~1_combout ),
	.sload(\MonDReg[8]~0_combout ),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_10),
	.prn(vcc));
defparam \MonDReg[10] .is_wysiwyg = "true";
defparam \MonDReg[10] .power_up = "low";

dffeas \MonDReg[9] (
	.clk(clk_clk),
	.d(jdo_12),
	.asdata(q_a_9),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[8]~1_combout ),
	.sload(\MonDReg[8]~0_combout ),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_9),
	.prn(vcc));
defparam \MonDReg[9] .is_wysiwyg = "true";
defparam \MonDReg[9] .power_up = "low";

dffeas \MonDReg[13] (
	.clk(clk_clk),
	.d(jdo_16),
	.asdata(q_a_13),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[8]~1_combout ),
	.sload(\MonDReg[8]~0_combout ),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_13),
	.prn(vcc));
defparam \MonDReg[13] .is_wysiwyg = "true";
defparam \MonDReg[13] .power_up = "low";

dffeas \MonDReg[14] (
	.clk(clk_clk),
	.d(jdo_17),
	.asdata(q_a_14),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[8]~1_combout ),
	.sload(\MonDReg[8]~0_combout ),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_14),
	.prn(vcc));
defparam \MonDReg[14] .is_wysiwyg = "true";
defparam \MonDReg[14] .power_up = "low";

dffeas waitrequest(
	.clk(clk_clk),
	.d(\waitrequest~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(waitrequest1),
	.prn(vcc));
defparam waitrequest.is_wysiwyg = "true";
defparam waitrequest.power_up = "low";

dffeas \MonDReg[0] (
	.clk(clk_clk),
	.d(\MonDReg~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_0),
	.prn(vcc));
defparam \MonDReg[0] .is_wysiwyg = "true";
defparam \MonDReg[0] .power_up = "low";

dffeas \MonDReg[1] (
	.clk(clk_clk),
	.d(\MonDReg~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_1),
	.prn(vcc));
defparam \MonDReg[1] .is_wysiwyg = "true";
defparam \MonDReg[1] .power_up = "low";

dffeas \MonDReg[3] (
	.clk(clk_clk),
	.d(\MonDReg~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_3),
	.prn(vcc));
defparam \MonDReg[3] .is_wysiwyg = "true";
defparam \MonDReg[3] .power_up = "low";

dffeas \MonDReg[18] (
	.clk(clk_clk),
	.d(\MonDReg~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_18),
	.prn(vcc));
defparam \MonDReg[18] .is_wysiwyg = "true";
defparam \MonDReg[18] .power_up = "low";

dffeas \MonDReg[4] (
	.clk(clk_clk),
	.d(\MonDReg~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_4),
	.prn(vcc));
defparam \MonDReg[4] .is_wysiwyg = "true";
defparam \MonDReg[4] .power_up = "low";

dffeas \MonDReg[22] (
	.clk(clk_clk),
	.d(\MonDReg~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_22),
	.prn(vcc));
defparam \MonDReg[22] .is_wysiwyg = "true";
defparam \MonDReg[22] .power_up = "low";

dffeas \MonDReg[5] (
	.clk(clk_clk),
	.d(\MonDReg~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_5),
	.prn(vcc));
defparam \MonDReg[5] .is_wysiwyg = "true";
defparam \MonDReg[5] .power_up = "low";

dffeas \MonDReg[29] (
	.clk(clk_clk),
	.d(\MonDReg~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_29),
	.prn(vcc));
defparam \MonDReg[29] .is_wysiwyg = "true";
defparam \MonDReg[29] .power_up = "low";

dffeas \MonDReg[8] (
	.clk(clk_clk),
	.d(\MonDReg~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_8),
	.prn(vcc));
defparam \MonDReg[8] .is_wysiwyg = "true";
defparam \MonDReg[8] .power_up = "low";

dffeas \MonDReg[15] (
	.clk(clk_clk),
	.d(\MonDReg~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!take_no_action_ocimem_a),
	.q(MonDReg_15),
	.prn(vcc));
defparam \MonDReg[15] .is_wysiwyg = "true";
defparam \MonDReg[15] .power_up = "low";

dffeas \MonDReg[12] (
	.clk(clk_clk),
	.d(\MonDReg~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_12),
	.prn(vcc));
defparam \MonDReg[12] .is_wysiwyg = "true";
defparam \MonDReg[12] .power_up = "low";

cyclonev_lcell_comb \Add0~1_wirecell (
	.dataa(!\Add0~1_sumout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~1_wirecell_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~1_wirecell .extended_lut = "off";
defparam \Add0~1_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \Add0~1_wirecell .shared_arith = "off";

dffeas \MonAReg[10] (
	.clk(clk_clk),
	.d(\Add0~1_wirecell_combout ),
	.asdata(jdo_17),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_a1),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[10]~q ),
	.prn(vcc));
defparam \MonAReg[10] .is_wysiwyg = "true";
defparam \MonAReg[10] .power_up = "low";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\MonAReg[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h00000000000000FF;
defparam \Add0~5 .shared_arith = "off";

dffeas \MonAReg[2] (
	.clk(clk_clk),
	.d(\Add0~5_sumout ),
	.asdata(jdo_26),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_a1),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[2]~q ),
	.prn(vcc));
defparam \MonAReg[2] .is_wysiwyg = "true";
defparam \MonAReg[2] .power_up = "low";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\MonAReg[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h00000000000000FF;
defparam \Add0~9 .shared_arith = "off";

dffeas \MonAReg[3] (
	.clk(clk_clk),
	.d(\Add0~9_sumout ),
	.asdata(jdo_27),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_a1),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[3]~q ),
	.prn(vcc));
defparam \MonAReg[3] .is_wysiwyg = "true";
defparam \MonAReg[3] .power_up = "low";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\MonAReg[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h00000000000000FF;
defparam \Add0~13 .shared_arith = "off";

dffeas \MonAReg[4] (
	.clk(clk_clk),
	.d(\Add0~13_sumout ),
	.asdata(jdo_28),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_a1),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[4]~q ),
	.prn(vcc));
defparam \MonAReg[4] .is_wysiwyg = "true";
defparam \MonAReg[4] .power_up = "low";

cyclonev_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\MonAReg[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h00000000000000FF;
defparam \Add0~21 .shared_arith = "off";

dffeas \MonAReg[5] (
	.clk(clk_clk),
	.d(\Add0~21_sumout ),
	.asdata(jdo_29),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_a1),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[5]~q ),
	.prn(vcc));
defparam \MonAReg[5] .is_wysiwyg = "true";
defparam \MonAReg[5] .power_up = "low";

cyclonev_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\MonAReg[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h00000000000000FF;
defparam \Add0~25 .shared_arith = "off";

dffeas \MonAReg[6] (
	.clk(clk_clk),
	.d(\Add0~25_sumout ),
	.asdata(jdo_30),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_a1),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[6]~q ),
	.prn(vcc));
defparam \MonAReg[6] .is_wysiwyg = "true";
defparam \MonAReg[6] .power_up = "low";

cyclonev_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\MonAReg[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout());
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h00000000000000FF;
defparam \Add0~29 .shared_arith = "off";

dffeas \MonAReg[7] (
	.clk(clk_clk),
	.d(\Add0~29_sumout ),
	.asdata(jdo_31),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_a1),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[7]~q ),
	.prn(vcc));
defparam \MonAReg[7] .is_wysiwyg = "true";
defparam \MonAReg[7] .power_up = "low";

cyclonev_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\MonAReg[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout());
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h00000000000000FF;
defparam \Add0~33 .shared_arith = "off";

dffeas \MonAReg[8] (
	.clk(clk_clk),
	.d(\Add0~33_sumout ),
	.asdata(jdo_32),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_a1),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[8]~q ),
	.prn(vcc));
defparam \MonAReg[8] .is_wysiwyg = "true";
defparam \MonAReg[8] .power_up = "low";

cyclonev_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\MonAReg[9]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h00000000000000FF;
defparam \Add0~17 .shared_arith = "off";

dffeas \MonAReg[9] (
	.clk(clk_clk),
	.d(\Add0~17_sumout ),
	.asdata(jdo_33),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_a1),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[9]~q ),
	.prn(vcc));
defparam \MonAReg[9] .is_wysiwyg = "true";
defparam \MonAReg[9] .power_up = "low";

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\MonAReg[10]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h00000000000000FF;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \jtag_ram_rd~0 (
	.dataa(!jdo_34),
	.datab(!take_no_action_ocimem_a),
	.datac(!jdo_17),
	.datad(!\Add0~1_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\jtag_ram_rd~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \jtag_ram_rd~0 .extended_lut = "off";
defparam \jtag_ram_rd~0 .lut_mask = 64'hB1FFB1FFB1FFB1FF;
defparam \jtag_ram_rd~0 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg[8]~0 (
	.dataa(!jdo_35),
	.datab(!take_action_ocimem_a),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg[8]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg[8]~0 .extended_lut = "off";
defparam \MonDReg[8]~0 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \MonDReg[8]~0 .shared_arith = "off";

dffeas jtag_ram_rd(
	.clk(clk_clk),
	.d(\jtag_ram_rd~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[8]~0_combout ),
	.q(\jtag_ram_rd~q ),
	.prn(vcc));
defparam jtag_ram_rd.is_wysiwyg = "true";
defparam jtag_ram_rd.power_up = "low";

dffeas jtag_ram_rd_d1(
	.clk(clk_clk),
	.d(\jtag_ram_rd~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jtag_ram_rd_d1~q ),
	.prn(vcc));
defparam jtag_ram_rd_d1.is_wysiwyg = "true";
defparam jtag_ram_rd_d1.power_up = "low";

cyclonev_lcell_comb \MonDReg[8]~1 (
	.dataa(!\jtag_ram_rd_d1~q ),
	.datab(!\MonDReg[8]~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg[8]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg[8]~1 .extended_lut = "off";
defparam \MonDReg[8]~1 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \MonDReg[8]~1 .shared_arith = "off";

dffeas jtag_rd(
	.clk(clk_clk),
	.d(take_no_action_ocimem_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[8]~0_combout ),
	.q(\jtag_rd~q ),
	.prn(vcc));
defparam jtag_rd.is_wysiwyg = "true";
defparam jtag_rd.power_up = "low";

dffeas jtag_rd_d1(
	.clk(clk_clk),
	.d(\jtag_rd~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jtag_rd_d1~q ),
	.prn(vcc));
defparam jtag_rd_d1.is_wysiwyg = "true";
defparam jtag_rd_d1.power_up = "low";

cyclonev_lcell_comb \MonDReg[0]~2 (
	.dataa(!jdo_35),
	.datab(!take_action_ocimem_a),
	.datac(!\jtag_rd_d1~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg[0]~2 .extended_lut = "off";
defparam \MonDReg[0]~2 .lut_mask = 64'h4747474747474747;
defparam \MonDReg[0]~2 .shared_arith = "off";

cyclonev_lcell_comb \jtag_ram_access~0 (
	.dataa(!jdo_34),
	.datab(!jdo_35),
	.datac(!take_action_ocimem_a),
	.datad(!jdo_17),
	.datae(!\Add0~1_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\jtag_ram_access~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \jtag_ram_access~0 .extended_lut = "off";
defparam \jtag_ram_access~0 .lut_mask = 64'hFF6FFFFFFF6FFFFF;
defparam \jtag_ram_access~0 .shared_arith = "off";

dffeas jtag_ram_access(
	.clk(clk_clk),
	.d(\jtag_ram_access~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jtag_ram_access~q ),
	.prn(vcc));
defparam jtag_ram_access.is_wysiwyg = "true";
defparam jtag_ram_access.power_up = "low";

cyclonev_lcell_comb \waitrequest~0 (
	.dataa(!address_8),
	.datab(!\jtag_ram_access~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\waitrequest~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \waitrequest~0 .extended_lut = "off";
defparam \waitrequest~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \waitrequest~0 .shared_arith = "off";

cyclonev_lcell_comb \avalon_ociram_readdata_ready~0 (
	.dataa(!waitrequest1),
	.datab(!write),
	.datac(!\waitrequest~0_combout ),
	.datad(!read),
	.datae(!\avalon_ociram_readdata_ready~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\avalon_ociram_readdata_ready~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \avalon_ociram_readdata_ready~0 .extended_lut = "off";
defparam \avalon_ociram_readdata_ready~0 .lut_mask = 64'hD1FFFFFFD1FFFFFF;
defparam \avalon_ociram_readdata_ready~0 .shared_arith = "off";

dffeas avalon_ociram_readdata_ready(
	.clk(clk_clk),
	.d(\avalon_ociram_readdata_ready~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\avalon_ociram_readdata_ready~q ),
	.prn(vcc));
defparam avalon_ociram_readdata_ready.is_wysiwyg = "true";
defparam avalon_ociram_readdata_ready.power_up = "low";

cyclonev_lcell_comb \waitrequest~1 (
	.dataa(!waitrequest1),
	.datab(!write),
	.datac(!\waitrequest~0_combout ),
	.datad(!read),
	.datae(!\avalon_ociram_readdata_ready~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\waitrequest~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \waitrequest~1 .extended_lut = "off";
defparam \waitrequest~1 .lut_mask = 64'hFFFFBF8FFFFFBF8F;
defparam \waitrequest~1 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg~16 (
	.dataa(!\MonAReg[4]~q ),
	.datab(!\MonAReg[3]~q ),
	.datac(!\jtag_ram_rd_d1~q ),
	.datad(!\MonAReg[2]~q ),
	.datae(!\MonDReg[8]~0_combout ),
	.dataf(!q_a_0),
	.datag(!jdo_3),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg~16 .extended_lut = "on";
defparam \MonDReg~16 .lut_mask = 64'hF7FBB77BF7FBB77B;
defparam \MonDReg~16 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~0 (
	.dataa(!\MonAReg[2]~q ),
	.datab(!\MonAReg[3]~q ),
	.datac(!\MonAReg[4]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~0 .extended_lut = "off";
defparam \Equal0~0 .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \Equal0~0 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg~3 (
	.dataa(!\jtag_ram_rd_d1~q ),
	.datab(!\MonDReg[8]~0_combout ),
	.datac(!\Equal0~0_combout ),
	.datad(!jdo_4),
	.datae(!q_a_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg~3 .extended_lut = "off";
defparam \MonDReg~3 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \MonDReg~3 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg~4 (
	.dataa(!\jtag_ram_rd_d1~q ),
	.datab(!\MonDReg[8]~0_combout ),
	.datac(!\Equal0~0_combout ),
	.datad(!jdo_6),
	.datae(!q_a_3),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg~4 .extended_lut = "off";
defparam \MonDReg~4 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \MonDReg~4 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg~5 (
	.dataa(!\MonAReg[2]~q ),
	.datab(!\MonAReg[3]~q ),
	.datac(!\MonAReg[4]~q ),
	.datad(!\jtag_ram_rd_d1~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg~5 .extended_lut = "off";
defparam \MonDReg~5 .lut_mask = 64'hFFFBFFFBFFFBFFFB;
defparam \MonDReg~5 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg~6 (
	.dataa(!jdo_21),
	.datab(!\jtag_ram_rd_d1~q ),
	.datac(!\MonDReg[8]~0_combout ),
	.datad(!q_a_18),
	.datae(!\MonDReg~5_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg~6 .extended_lut = "off";
defparam \MonDReg~6 .lut_mask = 64'h53FFFFFF53FFFFFF;
defparam \MonDReg~6 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg~7 (
	.dataa(!\MonAReg[2]~q ),
	.datab(!\MonAReg[3]~q ),
	.datac(!\MonAReg[4]~q ),
	.datad(!\jtag_ram_rd_d1~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg~7 .extended_lut = "off";
defparam \MonDReg~7 .lut_mask = 64'hFFFDFFFDFFFDFFFD;
defparam \MonDReg~7 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg~8 (
	.dataa(!\jtag_ram_rd_d1~q ),
	.datab(!\MonDReg[8]~0_combout ),
	.datac(!q_a_4),
	.datad(!jdo_7),
	.datae(!\MonDReg~7_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg~8 .extended_lut = "off";
defparam \MonDReg~8 .lut_mask = 64'h47FFFFFF47FFFFFF;
defparam \MonDReg~8 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg~9 (
	.dataa(!\jtag_ram_rd_d1~q ),
	.datab(!\MonDReg[8]~0_combout ),
	.datac(!jdo_25),
	.datad(!\MonDReg~5_combout ),
	.datae(!q_a_22),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg~9 .extended_lut = "off";
defparam \MonDReg~9 .lut_mask = 64'h47FFFFFF47FFFFFF;
defparam \MonDReg~9 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~1 (
	.dataa(!\MonAReg[2]~q ),
	.datab(!\MonAReg[3]~q ),
	.datac(!\MonAReg[4]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~1 .extended_lut = "off";
defparam \Equal0~1 .lut_mask = 64'hFEFEFEFEFEFEFEFE;
defparam \Equal0~1 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg~10 (
	.dataa(!\Equal0~1_combout ),
	.datab(!\jtag_ram_rd_d1~q ),
	.datac(!\MonDReg[8]~0_combout ),
	.datad(!q_a_5),
	.datae(!jdo_8),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg~10 .extended_lut = "off";
defparam \MonDReg~10 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \MonDReg~10 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg~11 (
	.dataa(!\jtag_ram_rd_d1~q ),
	.datab(!\MonDReg[8]~0_combout ),
	.datac(!\Equal0~0_combout ),
	.datad(!jdo_32),
	.datae(!q_a_29),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg~11 .extended_lut = "off";
defparam \MonDReg~11 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \MonDReg~11 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg~15 (
	.dataa(!\MonDReg[8]~0_combout ),
	.datab(!\jtag_ram_rd_d1~q ),
	.datac(!\MonAReg[4]~q ),
	.datad(!\MonAReg[2]~q ),
	.datae(!q_a_8),
	.dataf(!jdo_11),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg~15 .extended_lut = "off";
defparam \MonDReg~15 .lut_mask = 64'hF6FFFFFFFFFFFFFF;
defparam \MonDReg~15 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg~14 (
	.dataa(!\jtag_rd_d1~q ),
	.datab(!MonDReg_15),
	.datac(!\MonAReg[2]~q ),
	.datad(!\MonAReg[3]~q ),
	.datae(!\MonAReg[4]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg~14 .extended_lut = "off";
defparam \MonDReg~14 .lut_mask = 64'hFFB7FF7BFFB7FF7B;
defparam \MonDReg~14 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg~12 (
	.dataa(!\MonDReg[8]~0_combout ),
	.datab(!\jtag_rd_d1~q ),
	.datac(!jdo_18),
	.datad(!\jtag_ram_rd_d1~q ),
	.datae(!q_a_15),
	.dataf(!\MonDReg~14_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg~12 .extended_lut = "off";
defparam \MonDReg~12 .lut_mask = 64'h9F6FFFFFFFFFFFFF;
defparam \MonDReg~12 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg~13 (
	.dataa(!\jtag_ram_rd_d1~q ),
	.datab(!\MonDReg[8]~0_combout ),
	.datac(!\MonDReg~7_combout ),
	.datad(!q_a_12),
	.datae(!jdo_15),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg~13 .extended_lut = "off";
defparam \MonDReg~13 .lut_mask = 64'h47FFFFFF47FFFFFF;
defparam \MonDReg~13 .shared_arith = "off";

endmodule

module first_nios2_system_first_nios2_system_cpu_cpu_ociram_sp_ram_module (
	q_a_0,
	q_a_1,
	q_a_2,
	q_a_20,
	q_a_19,
	q_a_3,
	q_a_21,
	q_a_18,
	q_a_17,
	q_a_16,
	q_a_4,
	q_a_5,
	q_a_6,
	q_a_7,
	q_a_24,
	q_a_25,
	q_a_26,
	q_a_27,
	q_a_22,
	q_a_23,
	q_a_31,
	q_a_11,
	q_a_28,
	q_a_10,
	q_a_8,
	q_a_9,
	q_a_30,
	q_a_15,
	q_a_12,
	q_a_13,
	q_a_14,
	q_a_29,
	ociram_wr_en,
	ociram_reset_req,
	ociram_wr_data_0,
	ociram_addr_0,
	ociram_addr_1,
	ociram_addr_2,
	ociram_addr_3,
	ociram_addr_4,
	ociram_addr_5,
	ociram_addr_6,
	ociram_addr_7,
	ociram_byteenable_0,
	ociram_wr_data_1,
	ociram_wr_data_2,
	ociram_wr_data_20,
	ociram_byteenable_2,
	ociram_wr_data_19,
	ociram_wr_data_3,
	ociram_wr_data_21,
	ociram_wr_data_18,
	ociram_wr_data_17,
	ociram_wr_data_16,
	ociram_wr_data_4,
	ociram_wr_data_5,
	ociram_wr_data_6,
	ociram_wr_data_7,
	ociram_wr_data_24,
	ociram_byteenable_3,
	ociram_wr_data_25,
	ociram_wr_data_26,
	ociram_wr_data_27,
	ociram_wr_data_22,
	ociram_wr_data_23,
	ociram_wr_data_31,
	ociram_wr_data_11,
	ociram_byteenable_1,
	ociram_wr_data_28,
	ociram_wr_data_10,
	ociram_wr_data_8,
	ociram_wr_data_9,
	ociram_wr_data_30,
	ociram_wr_data_15,
	ociram_wr_data_12,
	ociram_wr_data_13,
	ociram_wr_data_14,
	ociram_wr_data_29,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	q_a_0;
output 	q_a_1;
output 	q_a_2;
output 	q_a_20;
output 	q_a_19;
output 	q_a_3;
output 	q_a_21;
output 	q_a_18;
output 	q_a_17;
output 	q_a_16;
output 	q_a_4;
output 	q_a_5;
output 	q_a_6;
output 	q_a_7;
output 	q_a_24;
output 	q_a_25;
output 	q_a_26;
output 	q_a_27;
output 	q_a_22;
output 	q_a_23;
output 	q_a_31;
output 	q_a_11;
output 	q_a_28;
output 	q_a_10;
output 	q_a_8;
output 	q_a_9;
output 	q_a_30;
output 	q_a_15;
output 	q_a_12;
output 	q_a_13;
output 	q_a_14;
output 	q_a_29;
input 	ociram_wr_en;
input 	ociram_reset_req;
input 	ociram_wr_data_0;
input 	ociram_addr_0;
input 	ociram_addr_1;
input 	ociram_addr_2;
input 	ociram_addr_3;
input 	ociram_addr_4;
input 	ociram_addr_5;
input 	ociram_addr_6;
input 	ociram_addr_7;
input 	ociram_byteenable_0;
input 	ociram_wr_data_1;
input 	ociram_wr_data_2;
input 	ociram_wr_data_20;
input 	ociram_byteenable_2;
input 	ociram_wr_data_19;
input 	ociram_wr_data_3;
input 	ociram_wr_data_21;
input 	ociram_wr_data_18;
input 	ociram_wr_data_17;
input 	ociram_wr_data_16;
input 	ociram_wr_data_4;
input 	ociram_wr_data_5;
input 	ociram_wr_data_6;
input 	ociram_wr_data_7;
input 	ociram_wr_data_24;
input 	ociram_byteenable_3;
input 	ociram_wr_data_25;
input 	ociram_wr_data_26;
input 	ociram_wr_data_27;
input 	ociram_wr_data_22;
input 	ociram_wr_data_23;
input 	ociram_wr_data_31;
input 	ociram_wr_data_11;
input 	ociram_byteenable_1;
input 	ociram_wr_data_28;
input 	ociram_wr_data_10;
input 	ociram_wr_data_8;
input 	ociram_wr_data_9;
input 	ociram_wr_data_30;
input 	ociram_wr_data_15;
input 	ociram_wr_data_12;
input 	ociram_wr_data_13;
input 	ociram_wr_data_14;
input 	ociram_wr_data_29;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



first_nios2_system_altsyncram_4 the_altsyncram(
	.q_a({q_a_31,q_a_30,q_a_29,q_a_28,q_a_27,q_a_26,q_a_25,q_a_24,q_a_23,q_a_22,q_a_21,q_a_20,q_a_19,q_a_18,q_a_17,q_a_16,q_a_15,q_a_14,q_a_13,q_a_12,q_a_11,q_a_10,q_a_9,q_a_8,q_a_7,q_a_6,q_a_5,q_a_4,q_a_3,q_a_2,q_a_1,q_a_0}),
	.wren_a(ociram_wr_en),
	.clocken0(ociram_reset_req),
	.data_a({ociram_wr_data_31,ociram_wr_data_30,ociram_wr_data_29,ociram_wr_data_28,ociram_wr_data_27,ociram_wr_data_26,ociram_wr_data_25,ociram_wr_data_24,ociram_wr_data_23,ociram_wr_data_22,ociram_wr_data_21,ociram_wr_data_20,ociram_wr_data_19,ociram_wr_data_18,ociram_wr_data_17,
ociram_wr_data_16,ociram_wr_data_15,ociram_wr_data_14,ociram_wr_data_13,ociram_wr_data_12,ociram_wr_data_11,ociram_wr_data_10,ociram_wr_data_9,ociram_wr_data_8,ociram_wr_data_7,ociram_wr_data_6,ociram_wr_data_5,ociram_wr_data_4,ociram_wr_data_3,ociram_wr_data_2,
ociram_wr_data_1,ociram_wr_data_0}),
	.address_a({gnd,gnd,gnd,gnd,gnd,ociram_addr_7,ociram_addr_6,ociram_addr_5,ociram_addr_4,ociram_addr_3,ociram_addr_2,ociram_addr_1,ociram_addr_0}),
	.byteena_a({ociram_byteenable_3,ociram_byteenable_2,ociram_byteenable_1,ociram_byteenable_0}),
	.clock0(clk_clk));

endmodule

module first_nios2_system_altsyncram_4 (
	q_a,
	wren_a,
	clocken0,
	data_a,
	address_a,
	byteena_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_a;
input 	wren_a;
input 	clocken0;
input 	[31:0] data_a;
input 	[12:0] address_a;
input 	[3:0] byteena_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



first_nios2_system_altsyncram_qid1 auto_generated(
	.q_a({q_a[31],q_a[30],q_a[29],q_a[28],q_a[27],q_a[26],q_a[25],q_a[24],q_a[23],q_a[22],q_a[21],q_a[20],q_a[19],q_a[18],q_a[17],q_a[16],q_a[15],q_a[14],q_a[13],q_a[12],q_a[11],q_a[10],q_a[9],q_a[8],q_a[7],q_a[6],q_a[5],q_a[4],q_a[3],q_a[2],q_a[1],q_a[0]}),
	.wren_a(wren_a),
	.clocken0(clocken0),
	.data_a({data_a[31],data_a[30],data_a[29],data_a[28],data_a[27],data_a[26],data_a[25],data_a[24],data_a[23],data_a[22],data_a[21],data_a[20],data_a[19],data_a[18],data_a[17],data_a[16],data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.address_a({address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.byteena_a({byteena_a[3],byteena_a[2],byteena_a[1],byteena_a[0]}),
	.clock0(clock0));

endmodule

module first_nios2_system_altsyncram_qid1 (
	q_a,
	wren_a,
	clocken0,
	data_a,
	address_a,
	byteena_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_a;
input 	wren_a;
input 	clocken0;
input 	[31:0] data_a;
input 	[7:0] address_a;
input 	[3:0] byteena_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTADATAOUT_bus;
wire [143:0] ram_block1a1_PORTADATAOUT_bus;
wire [143:0] ram_block1a2_PORTADATAOUT_bus;
wire [143:0] ram_block1a20_PORTADATAOUT_bus;
wire [143:0] ram_block1a19_PORTADATAOUT_bus;
wire [143:0] ram_block1a3_PORTADATAOUT_bus;
wire [143:0] ram_block1a21_PORTADATAOUT_bus;
wire [143:0] ram_block1a18_PORTADATAOUT_bus;
wire [143:0] ram_block1a17_PORTADATAOUT_bus;
wire [143:0] ram_block1a16_PORTADATAOUT_bus;
wire [143:0] ram_block1a4_PORTADATAOUT_bus;
wire [143:0] ram_block1a5_PORTADATAOUT_bus;
wire [143:0] ram_block1a6_PORTADATAOUT_bus;
wire [143:0] ram_block1a7_PORTADATAOUT_bus;
wire [143:0] ram_block1a24_PORTADATAOUT_bus;
wire [143:0] ram_block1a25_PORTADATAOUT_bus;
wire [143:0] ram_block1a26_PORTADATAOUT_bus;
wire [143:0] ram_block1a27_PORTADATAOUT_bus;
wire [143:0] ram_block1a22_PORTADATAOUT_bus;
wire [143:0] ram_block1a23_PORTADATAOUT_bus;
wire [143:0] ram_block1a31_PORTADATAOUT_bus;
wire [143:0] ram_block1a11_PORTADATAOUT_bus;
wire [143:0] ram_block1a28_PORTADATAOUT_bus;
wire [143:0] ram_block1a10_PORTADATAOUT_bus;
wire [143:0] ram_block1a8_PORTADATAOUT_bus;
wire [143:0] ram_block1a9_PORTADATAOUT_bus;
wire [143:0] ram_block1a30_PORTADATAOUT_bus;
wire [143:0] ram_block1a15_PORTADATAOUT_bus;
wire [143:0] ram_block1a12_PORTADATAOUT_bus;
wire [143:0] ram_block1a13_PORTADATAOUT_bus;
wire [143:0] ram_block1a14_PORTADATAOUT_bus;
wire [143:0] ram_block1a29_PORTADATAOUT_bus;

assign q_a[0] = ram_block1a0_PORTADATAOUT_bus[0];

assign q_a[1] = ram_block1a1_PORTADATAOUT_bus[0];

assign q_a[2] = ram_block1a2_PORTADATAOUT_bus[0];

assign q_a[20] = ram_block1a20_PORTADATAOUT_bus[0];

assign q_a[19] = ram_block1a19_PORTADATAOUT_bus[0];

assign q_a[3] = ram_block1a3_PORTADATAOUT_bus[0];

assign q_a[21] = ram_block1a21_PORTADATAOUT_bus[0];

assign q_a[18] = ram_block1a18_PORTADATAOUT_bus[0];

assign q_a[17] = ram_block1a17_PORTADATAOUT_bus[0];

assign q_a[16] = ram_block1a16_PORTADATAOUT_bus[0];

assign q_a[4] = ram_block1a4_PORTADATAOUT_bus[0];

assign q_a[5] = ram_block1a5_PORTADATAOUT_bus[0];

assign q_a[6] = ram_block1a6_PORTADATAOUT_bus[0];

assign q_a[7] = ram_block1a7_PORTADATAOUT_bus[0];

assign q_a[24] = ram_block1a24_PORTADATAOUT_bus[0];

assign q_a[25] = ram_block1a25_PORTADATAOUT_bus[0];

assign q_a[26] = ram_block1a26_PORTADATAOUT_bus[0];

assign q_a[27] = ram_block1a27_PORTADATAOUT_bus[0];

assign q_a[22] = ram_block1a22_PORTADATAOUT_bus[0];

assign q_a[23] = ram_block1a23_PORTADATAOUT_bus[0];

assign q_a[31] = ram_block1a31_PORTADATAOUT_bus[0];

assign q_a[11] = ram_block1a11_PORTADATAOUT_bus[0];

assign q_a[28] = ram_block1a28_PORTADATAOUT_bus[0];

assign q_a[10] = ram_block1a10_PORTADATAOUT_bus[0];

assign q_a[8] = ram_block1a8_PORTADATAOUT_bus[0];

assign q_a[9] = ram_block1a9_PORTADATAOUT_bus[0];

assign q_a[30] = ram_block1a30_PORTADATAOUT_bus[0];

assign q_a[15] = ram_block1a15_PORTADATAOUT_bus[0];

assign q_a[12] = ram_block1a12_PORTADATAOUT_bus[0];

assign q_a[13] = ram_block1a13_PORTADATAOUT_bus[0];

assign q_a[14] = ram_block1a14_PORTADATAOUT_bus[0];

assign q_a[29] = ram_block1a29_PORTADATAOUT_bus[0];

cyclonev_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a0_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_nios2_oci:the_first_nios2_system_cpu_cpu_nios2_oci|first_nios2_system_cpu_cpu_nios2_ocimem:the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram_module:first_nios2_system_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.operation_mode = "single_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 8;
defparam ram_block1a0.port_a_byte_enable_mask_width = 1;
defparam ram_block1a0.port_a_byte_size = 1;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 255;
defparam ram_block1a0.port_a_logical_ram_depth = 256;
defparam ram_block1a0.port_a_logical_ram_width = 32;
defparam ram_block1a0.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a0.ram_block_type = "auto";

cyclonev_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a1_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_nios2_oci:the_first_nios2_system_cpu_cpu_nios2_oci|first_nios2_system_cpu_cpu_nios2_ocimem:the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram_module:first_nios2_system_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.operation_mode = "single_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 8;
defparam ram_block1a1.port_a_byte_enable_mask_width = 1;
defparam ram_block1a1.port_a_byte_size = 1;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 255;
defparam ram_block1a1.port_a_logical_ram_depth = 256;
defparam ram_block1a1.port_a_logical_ram_width = 32;
defparam ram_block1a1.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a1.ram_block_type = "auto";

cyclonev_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a2_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_nios2_oci:the_first_nios2_system_cpu_cpu_nios2_oci|first_nios2_system_cpu_cpu_nios2_ocimem:the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram_module:first_nios2_system_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.operation_mode = "single_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 8;
defparam ram_block1a2.port_a_byte_enable_mask_width = 1;
defparam ram_block1a2.port_a_byte_size = 1;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 255;
defparam ram_block1a2.port_a_logical_ram_depth = 256;
defparam ram_block1a2.port_a_logical_ram_width = 32;
defparam ram_block1a2.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a2.ram_block_type = "auto";

cyclonev_ram_block ram_block1a20(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a20_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a20.clk0_core_clock_enable = "ena0";
defparam ram_block1a20.clk0_input_clock_enable = "ena0";
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_nios2_oci:the_first_nios2_system_cpu_cpu_nios2_oci|first_nios2_system_cpu_cpu_nios2_ocimem:the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram_module:first_nios2_system_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a20.operation_mode = "single_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 8;
defparam ram_block1a20.port_a_byte_enable_mask_width = 1;
defparam ram_block1a20.port_a_byte_size = 1;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 255;
defparam ram_block1a20.port_a_logical_ram_depth = 256;
defparam ram_block1a20.port_a_logical_ram_width = 32;
defparam ram_block1a20.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a20.ram_block_type = "auto";

cyclonev_ram_block ram_block1a19(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a19_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a19.clk0_core_clock_enable = "ena0";
defparam ram_block1a19.clk0_input_clock_enable = "ena0";
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_nios2_oci:the_first_nios2_system_cpu_cpu_nios2_oci|first_nios2_system_cpu_cpu_nios2_ocimem:the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram_module:first_nios2_system_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a19.operation_mode = "single_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 8;
defparam ram_block1a19.port_a_byte_enable_mask_width = 1;
defparam ram_block1a19.port_a_byte_size = 1;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 255;
defparam ram_block1a19.port_a_logical_ram_depth = 256;
defparam ram_block1a19.port_a_logical_ram_width = 32;
defparam ram_block1a19.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a19.ram_block_type = "auto";

cyclonev_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a3_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_nios2_oci:the_first_nios2_system_cpu_cpu_nios2_oci|first_nios2_system_cpu_cpu_nios2_ocimem:the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram_module:first_nios2_system_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.operation_mode = "single_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 8;
defparam ram_block1a3.port_a_byte_enable_mask_width = 1;
defparam ram_block1a3.port_a_byte_size = 1;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 255;
defparam ram_block1a3.port_a_logical_ram_depth = 256;
defparam ram_block1a3.port_a_logical_ram_width = 32;
defparam ram_block1a3.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a3.ram_block_type = "auto";

cyclonev_ram_block ram_block1a21(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a21_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a21.clk0_core_clock_enable = "ena0";
defparam ram_block1a21.clk0_input_clock_enable = "ena0";
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_nios2_oci:the_first_nios2_system_cpu_cpu_nios2_oci|first_nios2_system_cpu_cpu_nios2_ocimem:the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram_module:first_nios2_system_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a21.operation_mode = "single_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 8;
defparam ram_block1a21.port_a_byte_enable_mask_width = 1;
defparam ram_block1a21.port_a_byte_size = 1;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 255;
defparam ram_block1a21.port_a_logical_ram_depth = 256;
defparam ram_block1a21.port_a_logical_ram_width = 32;
defparam ram_block1a21.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a21.ram_block_type = "auto";

cyclonev_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a18_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a18.clk0_core_clock_enable = "ena0";
defparam ram_block1a18.clk0_input_clock_enable = "ena0";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_nios2_oci:the_first_nios2_system_cpu_cpu_nios2_oci|first_nios2_system_cpu_cpu_nios2_ocimem:the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram_module:first_nios2_system_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a18.operation_mode = "single_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 8;
defparam ram_block1a18.port_a_byte_enable_mask_width = 1;
defparam ram_block1a18.port_a_byte_size = 1;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 255;
defparam ram_block1a18.port_a_logical_ram_depth = 256;
defparam ram_block1a18.port_a_logical_ram_width = 32;
defparam ram_block1a18.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a18.ram_block_type = "auto";

cyclonev_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a17_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a17.clk0_core_clock_enable = "ena0";
defparam ram_block1a17.clk0_input_clock_enable = "ena0";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_nios2_oci:the_first_nios2_system_cpu_cpu_nios2_oci|first_nios2_system_cpu_cpu_nios2_ocimem:the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram_module:first_nios2_system_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a17.operation_mode = "single_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 8;
defparam ram_block1a17.port_a_byte_enable_mask_width = 1;
defparam ram_block1a17.port_a_byte_size = 1;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 255;
defparam ram_block1a17.port_a_logical_ram_depth = 256;
defparam ram_block1a17.port_a_logical_ram_width = 32;
defparam ram_block1a17.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a17.ram_block_type = "auto";

cyclonev_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a16_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a16.clk0_core_clock_enable = "ena0";
defparam ram_block1a16.clk0_input_clock_enable = "ena0";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_nios2_oci:the_first_nios2_system_cpu_cpu_nios2_oci|first_nios2_system_cpu_cpu_nios2_ocimem:the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram_module:first_nios2_system_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a16.operation_mode = "single_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 8;
defparam ram_block1a16.port_a_byte_enable_mask_width = 1;
defparam ram_block1a16.port_a_byte_size = 1;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 255;
defparam ram_block1a16.port_a_logical_ram_depth = 256;
defparam ram_block1a16.port_a_logical_ram_width = 32;
defparam ram_block1a16.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a16.ram_block_type = "auto";

cyclonev_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a4_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_nios2_oci:the_first_nios2_system_cpu_cpu_nios2_oci|first_nios2_system_cpu_cpu_nios2_ocimem:the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram_module:first_nios2_system_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.operation_mode = "single_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 8;
defparam ram_block1a4.port_a_byte_enable_mask_width = 1;
defparam ram_block1a4.port_a_byte_size = 1;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 255;
defparam ram_block1a4.port_a_logical_ram_depth = 256;
defparam ram_block1a4.port_a_logical_ram_width = 32;
defparam ram_block1a4.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a4.ram_block_type = "auto";

cyclonev_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a5_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_nios2_oci:the_first_nios2_system_cpu_cpu_nios2_oci|first_nios2_system_cpu_cpu_nios2_ocimem:the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram_module:first_nios2_system_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.operation_mode = "single_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 8;
defparam ram_block1a5.port_a_byte_enable_mask_width = 1;
defparam ram_block1a5.port_a_byte_size = 1;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 255;
defparam ram_block1a5.port_a_logical_ram_depth = 256;
defparam ram_block1a5.port_a_logical_ram_width = 32;
defparam ram_block1a5.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a5.ram_block_type = "auto";

cyclonev_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a6_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_nios2_oci:the_first_nios2_system_cpu_cpu_nios2_oci|first_nios2_system_cpu_cpu_nios2_ocimem:the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram_module:first_nios2_system_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.operation_mode = "single_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 8;
defparam ram_block1a6.port_a_byte_enable_mask_width = 1;
defparam ram_block1a6.port_a_byte_size = 1;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 255;
defparam ram_block1a6.port_a_logical_ram_depth = 256;
defparam ram_block1a6.port_a_logical_ram_width = 32;
defparam ram_block1a6.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a6.ram_block_type = "auto";

cyclonev_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a7_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_nios2_oci:the_first_nios2_system_cpu_cpu_nios2_oci|first_nios2_system_cpu_cpu_nios2_ocimem:the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram_module:first_nios2_system_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.operation_mode = "single_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 8;
defparam ram_block1a7.port_a_byte_enable_mask_width = 1;
defparam ram_block1a7.port_a_byte_size = 1;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 255;
defparam ram_block1a7.port_a_logical_ram_depth = 256;
defparam ram_block1a7.port_a_logical_ram_width = 32;
defparam ram_block1a7.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a7.ram_block_type = "auto";

cyclonev_ram_block ram_block1a24(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[24]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a24_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a24.clk0_core_clock_enable = "ena0";
defparam ram_block1a24.clk0_input_clock_enable = "ena0";
defparam ram_block1a24.data_interleave_offset_in_bits = 1;
defparam ram_block1a24.data_interleave_width_in_bits = 1;
defparam ram_block1a24.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_nios2_oci:the_first_nios2_system_cpu_cpu_nios2_oci|first_nios2_system_cpu_cpu_nios2_ocimem:the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram_module:first_nios2_system_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a24.operation_mode = "single_port";
defparam ram_block1a24.port_a_address_clear = "none";
defparam ram_block1a24.port_a_address_width = 8;
defparam ram_block1a24.port_a_byte_enable_mask_width = 1;
defparam ram_block1a24.port_a_byte_size = 1;
defparam ram_block1a24.port_a_data_out_clear = "none";
defparam ram_block1a24.port_a_data_out_clock = "none";
defparam ram_block1a24.port_a_data_width = 1;
defparam ram_block1a24.port_a_first_address = 0;
defparam ram_block1a24.port_a_first_bit_number = 24;
defparam ram_block1a24.port_a_last_address = 255;
defparam ram_block1a24.port_a_logical_ram_depth = 256;
defparam ram_block1a24.port_a_logical_ram_width = 32;
defparam ram_block1a24.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a24.ram_block_type = "auto";

cyclonev_ram_block ram_block1a25(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[25]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a25_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a25.clk0_core_clock_enable = "ena0";
defparam ram_block1a25.clk0_input_clock_enable = "ena0";
defparam ram_block1a25.data_interleave_offset_in_bits = 1;
defparam ram_block1a25.data_interleave_width_in_bits = 1;
defparam ram_block1a25.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_nios2_oci:the_first_nios2_system_cpu_cpu_nios2_oci|first_nios2_system_cpu_cpu_nios2_ocimem:the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram_module:first_nios2_system_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a25.operation_mode = "single_port";
defparam ram_block1a25.port_a_address_clear = "none";
defparam ram_block1a25.port_a_address_width = 8;
defparam ram_block1a25.port_a_byte_enable_mask_width = 1;
defparam ram_block1a25.port_a_byte_size = 1;
defparam ram_block1a25.port_a_data_out_clear = "none";
defparam ram_block1a25.port_a_data_out_clock = "none";
defparam ram_block1a25.port_a_data_width = 1;
defparam ram_block1a25.port_a_first_address = 0;
defparam ram_block1a25.port_a_first_bit_number = 25;
defparam ram_block1a25.port_a_last_address = 255;
defparam ram_block1a25.port_a_logical_ram_depth = 256;
defparam ram_block1a25.port_a_logical_ram_width = 32;
defparam ram_block1a25.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a25.ram_block_type = "auto";

cyclonev_ram_block ram_block1a26(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[26]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a26_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a26.clk0_core_clock_enable = "ena0";
defparam ram_block1a26.clk0_input_clock_enable = "ena0";
defparam ram_block1a26.data_interleave_offset_in_bits = 1;
defparam ram_block1a26.data_interleave_width_in_bits = 1;
defparam ram_block1a26.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_nios2_oci:the_first_nios2_system_cpu_cpu_nios2_oci|first_nios2_system_cpu_cpu_nios2_ocimem:the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram_module:first_nios2_system_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a26.operation_mode = "single_port";
defparam ram_block1a26.port_a_address_clear = "none";
defparam ram_block1a26.port_a_address_width = 8;
defparam ram_block1a26.port_a_byte_enable_mask_width = 1;
defparam ram_block1a26.port_a_byte_size = 1;
defparam ram_block1a26.port_a_data_out_clear = "none";
defparam ram_block1a26.port_a_data_out_clock = "none";
defparam ram_block1a26.port_a_data_width = 1;
defparam ram_block1a26.port_a_first_address = 0;
defparam ram_block1a26.port_a_first_bit_number = 26;
defparam ram_block1a26.port_a_last_address = 255;
defparam ram_block1a26.port_a_logical_ram_depth = 256;
defparam ram_block1a26.port_a_logical_ram_width = 32;
defparam ram_block1a26.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a26.ram_block_type = "auto";

cyclonev_ram_block ram_block1a27(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[27]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a27_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a27.clk0_core_clock_enable = "ena0";
defparam ram_block1a27.clk0_input_clock_enable = "ena0";
defparam ram_block1a27.data_interleave_offset_in_bits = 1;
defparam ram_block1a27.data_interleave_width_in_bits = 1;
defparam ram_block1a27.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_nios2_oci:the_first_nios2_system_cpu_cpu_nios2_oci|first_nios2_system_cpu_cpu_nios2_ocimem:the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram_module:first_nios2_system_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a27.operation_mode = "single_port";
defparam ram_block1a27.port_a_address_clear = "none";
defparam ram_block1a27.port_a_address_width = 8;
defparam ram_block1a27.port_a_byte_enable_mask_width = 1;
defparam ram_block1a27.port_a_byte_size = 1;
defparam ram_block1a27.port_a_data_out_clear = "none";
defparam ram_block1a27.port_a_data_out_clock = "none";
defparam ram_block1a27.port_a_data_width = 1;
defparam ram_block1a27.port_a_first_address = 0;
defparam ram_block1a27.port_a_first_bit_number = 27;
defparam ram_block1a27.port_a_last_address = 255;
defparam ram_block1a27.port_a_logical_ram_depth = 256;
defparam ram_block1a27.port_a_logical_ram_width = 32;
defparam ram_block1a27.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a27.ram_block_type = "auto";

cyclonev_ram_block ram_block1a22(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[22]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a22_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a22.clk0_core_clock_enable = "ena0";
defparam ram_block1a22.clk0_input_clock_enable = "ena0";
defparam ram_block1a22.data_interleave_offset_in_bits = 1;
defparam ram_block1a22.data_interleave_width_in_bits = 1;
defparam ram_block1a22.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_nios2_oci:the_first_nios2_system_cpu_cpu_nios2_oci|first_nios2_system_cpu_cpu_nios2_ocimem:the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram_module:first_nios2_system_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a22.operation_mode = "single_port";
defparam ram_block1a22.port_a_address_clear = "none";
defparam ram_block1a22.port_a_address_width = 8;
defparam ram_block1a22.port_a_byte_enable_mask_width = 1;
defparam ram_block1a22.port_a_byte_size = 1;
defparam ram_block1a22.port_a_data_out_clear = "none";
defparam ram_block1a22.port_a_data_out_clock = "none";
defparam ram_block1a22.port_a_data_width = 1;
defparam ram_block1a22.port_a_first_address = 0;
defparam ram_block1a22.port_a_first_bit_number = 22;
defparam ram_block1a22.port_a_last_address = 255;
defparam ram_block1a22.port_a_logical_ram_depth = 256;
defparam ram_block1a22.port_a_logical_ram_width = 32;
defparam ram_block1a22.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a22.ram_block_type = "auto";

cyclonev_ram_block ram_block1a23(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[23]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a23_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a23.clk0_core_clock_enable = "ena0";
defparam ram_block1a23.clk0_input_clock_enable = "ena0";
defparam ram_block1a23.data_interleave_offset_in_bits = 1;
defparam ram_block1a23.data_interleave_width_in_bits = 1;
defparam ram_block1a23.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_nios2_oci:the_first_nios2_system_cpu_cpu_nios2_oci|first_nios2_system_cpu_cpu_nios2_ocimem:the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram_module:first_nios2_system_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a23.operation_mode = "single_port";
defparam ram_block1a23.port_a_address_clear = "none";
defparam ram_block1a23.port_a_address_width = 8;
defparam ram_block1a23.port_a_byte_enable_mask_width = 1;
defparam ram_block1a23.port_a_byte_size = 1;
defparam ram_block1a23.port_a_data_out_clear = "none";
defparam ram_block1a23.port_a_data_out_clock = "none";
defparam ram_block1a23.port_a_data_width = 1;
defparam ram_block1a23.port_a_first_address = 0;
defparam ram_block1a23.port_a_first_bit_number = 23;
defparam ram_block1a23.port_a_last_address = 255;
defparam ram_block1a23.port_a_logical_ram_depth = 256;
defparam ram_block1a23.port_a_logical_ram_width = 32;
defparam ram_block1a23.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a23.ram_block_type = "auto";

cyclonev_ram_block ram_block1a31(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a31_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a31.clk0_core_clock_enable = "ena0";
defparam ram_block1a31.clk0_input_clock_enable = "ena0";
defparam ram_block1a31.data_interleave_offset_in_bits = 1;
defparam ram_block1a31.data_interleave_width_in_bits = 1;
defparam ram_block1a31.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_nios2_oci:the_first_nios2_system_cpu_cpu_nios2_oci|first_nios2_system_cpu_cpu_nios2_ocimem:the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram_module:first_nios2_system_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a31.operation_mode = "single_port";
defparam ram_block1a31.port_a_address_clear = "none";
defparam ram_block1a31.port_a_address_width = 8;
defparam ram_block1a31.port_a_byte_enable_mask_width = 1;
defparam ram_block1a31.port_a_byte_size = 1;
defparam ram_block1a31.port_a_data_out_clear = "none";
defparam ram_block1a31.port_a_data_out_clock = "none";
defparam ram_block1a31.port_a_data_width = 1;
defparam ram_block1a31.port_a_first_address = 0;
defparam ram_block1a31.port_a_first_bit_number = 31;
defparam ram_block1a31.port_a_last_address = 255;
defparam ram_block1a31.port_a_logical_ram_depth = 256;
defparam ram_block1a31.port_a_logical_ram_width = 32;
defparam ram_block1a31.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a31.ram_block_type = "auto";

cyclonev_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a11_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.clk0_input_clock_enable = "ena0";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_nios2_oci:the_first_nios2_system_cpu_cpu_nios2_oci|first_nios2_system_cpu_cpu_nios2_ocimem:the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram_module:first_nios2_system_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.operation_mode = "single_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 8;
defparam ram_block1a11.port_a_byte_enable_mask_width = 1;
defparam ram_block1a11.port_a_byte_size = 1;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 255;
defparam ram_block1a11.port_a_logical_ram_depth = 256;
defparam ram_block1a11.port_a_logical_ram_width = 32;
defparam ram_block1a11.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a11.ram_block_type = "auto";

cyclonev_ram_block ram_block1a28(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[28]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a28_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a28.clk0_core_clock_enable = "ena0";
defparam ram_block1a28.clk0_input_clock_enable = "ena0";
defparam ram_block1a28.data_interleave_offset_in_bits = 1;
defparam ram_block1a28.data_interleave_width_in_bits = 1;
defparam ram_block1a28.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_nios2_oci:the_first_nios2_system_cpu_cpu_nios2_oci|first_nios2_system_cpu_cpu_nios2_ocimem:the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram_module:first_nios2_system_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a28.operation_mode = "single_port";
defparam ram_block1a28.port_a_address_clear = "none";
defparam ram_block1a28.port_a_address_width = 8;
defparam ram_block1a28.port_a_byte_enable_mask_width = 1;
defparam ram_block1a28.port_a_byte_size = 1;
defparam ram_block1a28.port_a_data_out_clear = "none";
defparam ram_block1a28.port_a_data_out_clock = "none";
defparam ram_block1a28.port_a_data_width = 1;
defparam ram_block1a28.port_a_first_address = 0;
defparam ram_block1a28.port_a_first_bit_number = 28;
defparam ram_block1a28.port_a_last_address = 255;
defparam ram_block1a28.port_a_logical_ram_depth = 256;
defparam ram_block1a28.port_a_logical_ram_width = 32;
defparam ram_block1a28.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a28.ram_block_type = "auto";

cyclonev_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a10_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.clk0_input_clock_enable = "ena0";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_nios2_oci:the_first_nios2_system_cpu_cpu_nios2_oci|first_nios2_system_cpu_cpu_nios2_ocimem:the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram_module:first_nios2_system_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.operation_mode = "single_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 8;
defparam ram_block1a10.port_a_byte_enable_mask_width = 1;
defparam ram_block1a10.port_a_byte_size = 1;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 255;
defparam ram_block1a10.port_a_logical_ram_depth = 256;
defparam ram_block1a10.port_a_logical_ram_width = 32;
defparam ram_block1a10.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a10.ram_block_type = "auto";

cyclonev_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a8_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk0_input_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_nios2_oci:the_first_nios2_system_cpu_cpu_nios2_oci|first_nios2_system_cpu_cpu_nios2_ocimem:the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram_module:first_nios2_system_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.operation_mode = "single_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 8;
defparam ram_block1a8.port_a_byte_enable_mask_width = 1;
defparam ram_block1a8.port_a_byte_size = 1;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 255;
defparam ram_block1a8.port_a_logical_ram_depth = 256;
defparam ram_block1a8.port_a_logical_ram_width = 32;
defparam ram_block1a8.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a8.ram_block_type = "auto";

cyclonev_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a9_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk0_input_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_nios2_oci:the_first_nios2_system_cpu_cpu_nios2_oci|first_nios2_system_cpu_cpu_nios2_ocimem:the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram_module:first_nios2_system_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.operation_mode = "single_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 8;
defparam ram_block1a9.port_a_byte_enable_mask_width = 1;
defparam ram_block1a9.port_a_byte_size = 1;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 255;
defparam ram_block1a9.port_a_logical_ram_depth = 256;
defparam ram_block1a9.port_a_logical_ram_width = 32;
defparam ram_block1a9.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a9.ram_block_type = "auto";

cyclonev_ram_block ram_block1a30(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[30]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a30_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a30.clk0_core_clock_enable = "ena0";
defparam ram_block1a30.clk0_input_clock_enable = "ena0";
defparam ram_block1a30.data_interleave_offset_in_bits = 1;
defparam ram_block1a30.data_interleave_width_in_bits = 1;
defparam ram_block1a30.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_nios2_oci:the_first_nios2_system_cpu_cpu_nios2_oci|first_nios2_system_cpu_cpu_nios2_ocimem:the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram_module:first_nios2_system_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a30.operation_mode = "single_port";
defparam ram_block1a30.port_a_address_clear = "none";
defparam ram_block1a30.port_a_address_width = 8;
defparam ram_block1a30.port_a_byte_enable_mask_width = 1;
defparam ram_block1a30.port_a_byte_size = 1;
defparam ram_block1a30.port_a_data_out_clear = "none";
defparam ram_block1a30.port_a_data_out_clock = "none";
defparam ram_block1a30.port_a_data_width = 1;
defparam ram_block1a30.port_a_first_address = 0;
defparam ram_block1a30.port_a_first_bit_number = 30;
defparam ram_block1a30.port_a_last_address = 255;
defparam ram_block1a30.port_a_logical_ram_depth = 256;
defparam ram_block1a30.port_a_logical_ram_width = 32;
defparam ram_block1a30.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a30.ram_block_type = "auto";

cyclonev_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a15_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.clk0_input_clock_enable = "ena0";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_nios2_oci:the_first_nios2_system_cpu_cpu_nios2_oci|first_nios2_system_cpu_cpu_nios2_ocimem:the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram_module:first_nios2_system_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.operation_mode = "single_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 8;
defparam ram_block1a15.port_a_byte_enable_mask_width = 1;
defparam ram_block1a15.port_a_byte_size = 1;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 255;
defparam ram_block1a15.port_a_logical_ram_depth = 256;
defparam ram_block1a15.port_a_logical_ram_width = 32;
defparam ram_block1a15.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a15.ram_block_type = "auto";

cyclonev_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a12_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.clk0_input_clock_enable = "ena0";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_nios2_oci:the_first_nios2_system_cpu_cpu_nios2_oci|first_nios2_system_cpu_cpu_nios2_ocimem:the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram_module:first_nios2_system_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.operation_mode = "single_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 8;
defparam ram_block1a12.port_a_byte_enable_mask_width = 1;
defparam ram_block1a12.port_a_byte_size = 1;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 255;
defparam ram_block1a12.port_a_logical_ram_depth = 256;
defparam ram_block1a12.port_a_logical_ram_width = 32;
defparam ram_block1a12.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a12.ram_block_type = "auto";

cyclonev_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a13_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.clk0_input_clock_enable = "ena0";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_nios2_oci:the_first_nios2_system_cpu_cpu_nios2_oci|first_nios2_system_cpu_cpu_nios2_ocimem:the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram_module:first_nios2_system_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.operation_mode = "single_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 8;
defparam ram_block1a13.port_a_byte_enable_mask_width = 1;
defparam ram_block1a13.port_a_byte_size = 1;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 255;
defparam ram_block1a13.port_a_logical_ram_depth = 256;
defparam ram_block1a13.port_a_logical_ram_width = 32;
defparam ram_block1a13.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a13.ram_block_type = "auto";

cyclonev_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a14_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.clk0_input_clock_enable = "ena0";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_nios2_oci:the_first_nios2_system_cpu_cpu_nios2_oci|first_nios2_system_cpu_cpu_nios2_ocimem:the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram_module:first_nios2_system_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.operation_mode = "single_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 8;
defparam ram_block1a14.port_a_byte_enable_mask_width = 1;
defparam ram_block1a14.port_a_byte_size = 1;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 255;
defparam ram_block1a14.port_a_logical_ram_depth = 256;
defparam ram_block1a14.port_a_logical_ram_width = 32;
defparam ram_block1a14.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a14.ram_block_type = "auto";

cyclonev_ram_block ram_block1a29(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[29]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a29_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a29.clk0_core_clock_enable = "ena0";
defparam ram_block1a29.clk0_input_clock_enable = "ena0";
defparam ram_block1a29.data_interleave_offset_in_bits = 1;
defparam ram_block1a29.data_interleave_width_in_bits = 1;
defparam ram_block1a29.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_nios2_oci:the_first_nios2_system_cpu_cpu_nios2_oci|first_nios2_system_cpu_cpu_nios2_ocimem:the_first_nios2_system_cpu_cpu_nios2_ocimem|first_nios2_system_cpu_cpu_ociram_sp_ram_module:first_nios2_system_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a29.operation_mode = "single_port";
defparam ram_block1a29.port_a_address_clear = "none";
defparam ram_block1a29.port_a_address_width = 8;
defparam ram_block1a29.port_a_byte_enable_mask_width = 1;
defparam ram_block1a29.port_a_byte_size = 1;
defparam ram_block1a29.port_a_data_out_clear = "none";
defparam ram_block1a29.port_a_data_out_clock = "none";
defparam ram_block1a29.port_a_data_width = 1;
defparam ram_block1a29.port_a_first_address = 0;
defparam ram_block1a29.port_a_first_bit_number = 29;
defparam ram_block1a29.port_a_last_address = 255;
defparam ram_block1a29.port_a_logical_ram_depth = 256;
defparam ram_block1a29.port_a_logical_ram_width = 32;
defparam ram_block1a29.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a29.ram_block_type = "auto";

endmodule

module first_nios2_system_first_nios2_system_cpu_cpu_register_bank_a_module (
	q_b_3,
	q_b_22,
	q_b_23,
	q_b_24,
	q_b_0,
	q_b_25,
	q_b_2,
	q_b_31,
	q_b_7,
	q_b_21,
	q_b_11,
	q_b_28,
	q_b_10,
	q_b_27,
	q_b_8,
	q_b_9,
	q_b_4,
	q_b_5,
	q_b_6,
	q_b_26,
	q_b_20,
	q_b_19,
	q_b_17,
	q_b_30,
	q_b_1,
	q_b_18,
	q_b_16,
	q_b_15,
	q_b_12,
	q_b_13,
	q_b_14,
	q_b_29,
	A_wr_data_unfiltered_0,
	A_wr_data_unfiltered_1,
	A_wr_data_unfiltered_2,
	A_wr_data_unfiltered_3,
	A_wr_data_unfiltered_4,
	A_wr_data_unfiltered_5,
	A_wr_data_unfiltered_6,
	A_wr_data_unfiltered_7,
	A_wr_data_unfiltered_22,
	A_wr_data_unfiltered_23,
	A_wr_data_unfiltered_24,
	A_wr_data_unfiltered_25,
	A_wr_data_unfiltered_31,
	A_wr_data_unfiltered_21,
	A_wr_data_unfiltered_11,
	A_wr_data_unfiltered_28,
	A_wr_data_unfiltered_10,
	A_wr_data_unfiltered_27,
	A_wr_data_unfiltered_8,
	A_wr_data_unfiltered_9,
	A_wr_data_unfiltered_26,
	A_wr_data_unfiltered_20,
	A_wr_data_unfiltered_19,
	A_wr_data_unfiltered_17,
	A_wr_data_unfiltered_30,
	A_wr_data_unfiltered_18,
	A_wr_data_unfiltered_16,
	A_wr_data_unfiltered_15,
	A_wr_data_unfiltered_12,
	A_wr_data_unfiltered_13,
	A_wr_data_unfiltered_14,
	A_wr_data_unfiltered_29,
	A_wr_dst_reg,
	A_dst_regnum,
	A_dst_regnum1,
	A_dst_regnum2,
	A_dst_regnum3,
	A_dst_regnum4,
	rf_a_rd_port_addr_0,
	rf_a_rd_port_addr_1,
	rf_a_rd_port_addr_2,
	rf_a_rd_port_addr_3,
	rf_a_rd_port_addr_4,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_3;
output 	q_b_22;
output 	q_b_23;
output 	q_b_24;
output 	q_b_0;
output 	q_b_25;
output 	q_b_2;
output 	q_b_31;
output 	q_b_7;
output 	q_b_21;
output 	q_b_11;
output 	q_b_28;
output 	q_b_10;
output 	q_b_27;
output 	q_b_8;
output 	q_b_9;
output 	q_b_4;
output 	q_b_5;
output 	q_b_6;
output 	q_b_26;
output 	q_b_20;
output 	q_b_19;
output 	q_b_17;
output 	q_b_30;
output 	q_b_1;
output 	q_b_18;
output 	q_b_16;
output 	q_b_15;
output 	q_b_12;
output 	q_b_13;
output 	q_b_14;
output 	q_b_29;
input 	A_wr_data_unfiltered_0;
input 	A_wr_data_unfiltered_1;
input 	A_wr_data_unfiltered_2;
input 	A_wr_data_unfiltered_3;
input 	A_wr_data_unfiltered_4;
input 	A_wr_data_unfiltered_5;
input 	A_wr_data_unfiltered_6;
input 	A_wr_data_unfiltered_7;
input 	A_wr_data_unfiltered_22;
input 	A_wr_data_unfiltered_23;
input 	A_wr_data_unfiltered_24;
input 	A_wr_data_unfiltered_25;
input 	A_wr_data_unfiltered_31;
input 	A_wr_data_unfiltered_21;
input 	A_wr_data_unfiltered_11;
input 	A_wr_data_unfiltered_28;
input 	A_wr_data_unfiltered_10;
input 	A_wr_data_unfiltered_27;
input 	A_wr_data_unfiltered_8;
input 	A_wr_data_unfiltered_9;
input 	A_wr_data_unfiltered_26;
input 	A_wr_data_unfiltered_20;
input 	A_wr_data_unfiltered_19;
input 	A_wr_data_unfiltered_17;
input 	A_wr_data_unfiltered_30;
input 	A_wr_data_unfiltered_18;
input 	A_wr_data_unfiltered_16;
input 	A_wr_data_unfiltered_15;
input 	A_wr_data_unfiltered_12;
input 	A_wr_data_unfiltered_13;
input 	A_wr_data_unfiltered_14;
input 	A_wr_data_unfiltered_29;
input 	A_wr_dst_reg;
input 	A_dst_regnum;
input 	A_dst_regnum1;
input 	A_dst_regnum2;
input 	A_dst_regnum3;
input 	A_dst_regnum4;
input 	rf_a_rd_port_addr_0;
input 	rf_a_rd_port_addr_1;
input 	rf_a_rd_port_addr_2;
input 	rf_a_rd_port_addr_3;
input 	rf_a_rd_port_addr_4;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



first_nios2_system_altsyncram_5 the_altsyncram(
	.q_b({q_b_31,q_b_30,q_b_29,q_b_28,q_b_27,q_b_26,q_b_25,q_b_24,q_b_23,q_b_22,q_b_21,q_b_20,q_b_19,q_b_18,q_b_17,q_b_16,q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.data_a({A_wr_data_unfiltered_31,A_wr_data_unfiltered_30,A_wr_data_unfiltered_29,A_wr_data_unfiltered_28,A_wr_data_unfiltered_27,A_wr_data_unfiltered_26,A_wr_data_unfiltered_25,A_wr_data_unfiltered_24,A_wr_data_unfiltered_23,A_wr_data_unfiltered_22,A_wr_data_unfiltered_21,
A_wr_data_unfiltered_20,A_wr_data_unfiltered_19,A_wr_data_unfiltered_18,A_wr_data_unfiltered_17,A_wr_data_unfiltered_16,A_wr_data_unfiltered_15,A_wr_data_unfiltered_14,A_wr_data_unfiltered_13,A_wr_data_unfiltered_12,A_wr_data_unfiltered_11,A_wr_data_unfiltered_10,
A_wr_data_unfiltered_9,A_wr_data_unfiltered_8,A_wr_data_unfiltered_7,A_wr_data_unfiltered_6,A_wr_data_unfiltered_5,A_wr_data_unfiltered_4,A_wr_data_unfiltered_3,A_wr_data_unfiltered_2,A_wr_data_unfiltered_1,A_wr_data_unfiltered_0}),
	.wren_a(A_wr_dst_reg),
	.address_a({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,A_dst_regnum4,A_dst_regnum3,A_dst_regnum2,A_dst_regnum1,A_dst_regnum}),
	.address_b({gnd,gnd,gnd,gnd,rf_a_rd_port_addr_4,rf_a_rd_port_addr_3,rf_a_rd_port_addr_2,rf_a_rd_port_addr_1,rf_a_rd_port_addr_0}),
	.clock0(clk_clk));

endmodule

module first_nios2_system_altsyncram_5 (
	q_b,
	data_a,
	wren_a,
	address_a,
	address_b,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_b;
input 	[31:0] data_a;
input 	wren_a;
input 	[12:0] address_a;
input 	[8:0] address_b;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



first_nios2_system_altsyncram_voi1 auto_generated(
	.q_b({q_b[31],q_b[30],q_b[29],q_b[28],q_b[27],q_b[26],q_b[25],q_b[24],q_b[23],q_b[22],q_b[21],q_b[20],q_b[19],q_b[18],q_b[17],q_b[16],q_b[15],q_b[14],q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.data_a({data_a[31],data_a[30],data_a[29],data_a[28],data_a[27],data_a[26],data_a[25],data_a[24],data_a[23],data_a[22],data_a[21],data_a[20],data_a[19],data_a[18],data_a[17],data_a[16],data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.wren_a(wren_a),
	.address_a({address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.address_b({address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.clock0(clock0));

endmodule

module first_nios2_system_altsyncram_voi1 (
	q_b,
	data_a,
	wren_a,
	address_a,
	address_b,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_b;
input 	[31:0] data_a;
input 	wren_a;
input 	[4:0] address_a;
input 	[4:0] address_b;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a22_PORTBDATAOUT_bus;
wire [143:0] ram_block1a23_PORTBDATAOUT_bus;
wire [143:0] ram_block1a24_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a25_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a31_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a21_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a28_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a27_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a26_PORTBDATAOUT_bus;
wire [143:0] ram_block1a20_PORTBDATAOUT_bus;
wire [143:0] ram_block1a19_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;
wire [143:0] ram_block1a30_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a29_PORTBDATAOUT_bus;

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[22] = ram_block1a22_PORTBDATAOUT_bus[0];

assign q_b[23] = ram_block1a23_PORTBDATAOUT_bus[0];

assign q_b[24] = ram_block1a24_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[25] = ram_block1a25_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[31] = ram_block1a31_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[21] = ram_block1a21_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[28] = ram_block1a28_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[27] = ram_block1a27_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[26] = ram_block1a26_PORTBDATAOUT_bus[0];

assign q_b[20] = ram_block1a20_PORTBDATAOUT_bus[0];

assign q_b[19] = ram_block1a19_PORTBDATAOUT_bus[0];

assign q_b[17] = ram_block1a17_PORTBDATAOUT_bus[0];

assign q_b[30] = ram_block1a30_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[18] = ram_block1a18_PORTBDATAOUT_bus[0];

assign q_b[16] = ram_block1a16_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[29] = ram_block1a29_PORTBDATAOUT_bus[0];

cyclonev_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_register_bank_a_module:first_nios2_system_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_voi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "old";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 5;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 31;
defparam ram_block1a3.port_a_logical_ram_depth = 32;
defparam ram_block1a3.port_a_logical_ram_width = 32;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock0";
defparam ram_block1a3.port_b_address_width = 5;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "none";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 31;
defparam ram_block1a3.port_b_logical_ram_depth = 32;
defparam ram_block1a3.port_b_logical_ram_width = 32;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock0";
defparam ram_block1a3.ram_block_type = "auto";

cyclonev_ram_block ram_block1a22(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[22]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a22_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a22.data_interleave_offset_in_bits = 1;
defparam ram_block1a22.data_interleave_width_in_bits = 1;
defparam ram_block1a22.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_register_bank_a_module:first_nios2_system_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_voi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a22.mixed_port_feed_through_mode = "old";
defparam ram_block1a22.operation_mode = "dual_port";
defparam ram_block1a22.port_a_address_clear = "none";
defparam ram_block1a22.port_a_address_width = 5;
defparam ram_block1a22.port_a_data_out_clear = "none";
defparam ram_block1a22.port_a_data_out_clock = "none";
defparam ram_block1a22.port_a_data_width = 1;
defparam ram_block1a22.port_a_first_address = 0;
defparam ram_block1a22.port_a_first_bit_number = 22;
defparam ram_block1a22.port_a_last_address = 31;
defparam ram_block1a22.port_a_logical_ram_depth = 32;
defparam ram_block1a22.port_a_logical_ram_width = 32;
defparam ram_block1a22.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a22.port_b_address_clear = "none";
defparam ram_block1a22.port_b_address_clock = "clock0";
defparam ram_block1a22.port_b_address_width = 5;
defparam ram_block1a22.port_b_data_out_clear = "none";
defparam ram_block1a22.port_b_data_out_clock = "none";
defparam ram_block1a22.port_b_data_width = 1;
defparam ram_block1a22.port_b_first_address = 0;
defparam ram_block1a22.port_b_first_bit_number = 22;
defparam ram_block1a22.port_b_last_address = 31;
defparam ram_block1a22.port_b_logical_ram_depth = 32;
defparam ram_block1a22.port_b_logical_ram_width = 32;
defparam ram_block1a22.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a22.port_b_read_enable_clock = "clock0";
defparam ram_block1a22.ram_block_type = "auto";

cyclonev_ram_block ram_block1a23(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[23]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a23_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a23.data_interleave_offset_in_bits = 1;
defparam ram_block1a23.data_interleave_width_in_bits = 1;
defparam ram_block1a23.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_register_bank_a_module:first_nios2_system_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_voi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a23.mixed_port_feed_through_mode = "old";
defparam ram_block1a23.operation_mode = "dual_port";
defparam ram_block1a23.port_a_address_clear = "none";
defparam ram_block1a23.port_a_address_width = 5;
defparam ram_block1a23.port_a_data_out_clear = "none";
defparam ram_block1a23.port_a_data_out_clock = "none";
defparam ram_block1a23.port_a_data_width = 1;
defparam ram_block1a23.port_a_first_address = 0;
defparam ram_block1a23.port_a_first_bit_number = 23;
defparam ram_block1a23.port_a_last_address = 31;
defparam ram_block1a23.port_a_logical_ram_depth = 32;
defparam ram_block1a23.port_a_logical_ram_width = 32;
defparam ram_block1a23.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a23.port_b_address_clear = "none";
defparam ram_block1a23.port_b_address_clock = "clock0";
defparam ram_block1a23.port_b_address_width = 5;
defparam ram_block1a23.port_b_data_out_clear = "none";
defparam ram_block1a23.port_b_data_out_clock = "none";
defparam ram_block1a23.port_b_data_width = 1;
defparam ram_block1a23.port_b_first_address = 0;
defparam ram_block1a23.port_b_first_bit_number = 23;
defparam ram_block1a23.port_b_last_address = 31;
defparam ram_block1a23.port_b_logical_ram_depth = 32;
defparam ram_block1a23.port_b_logical_ram_width = 32;
defparam ram_block1a23.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a23.port_b_read_enable_clock = "clock0";
defparam ram_block1a23.ram_block_type = "auto";

cyclonev_ram_block ram_block1a24(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[24]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a24_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a24.data_interleave_offset_in_bits = 1;
defparam ram_block1a24.data_interleave_width_in_bits = 1;
defparam ram_block1a24.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_register_bank_a_module:first_nios2_system_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_voi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a24.mixed_port_feed_through_mode = "old";
defparam ram_block1a24.operation_mode = "dual_port";
defparam ram_block1a24.port_a_address_clear = "none";
defparam ram_block1a24.port_a_address_width = 5;
defparam ram_block1a24.port_a_data_out_clear = "none";
defparam ram_block1a24.port_a_data_out_clock = "none";
defparam ram_block1a24.port_a_data_width = 1;
defparam ram_block1a24.port_a_first_address = 0;
defparam ram_block1a24.port_a_first_bit_number = 24;
defparam ram_block1a24.port_a_last_address = 31;
defparam ram_block1a24.port_a_logical_ram_depth = 32;
defparam ram_block1a24.port_a_logical_ram_width = 32;
defparam ram_block1a24.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a24.port_b_address_clear = "none";
defparam ram_block1a24.port_b_address_clock = "clock0";
defparam ram_block1a24.port_b_address_width = 5;
defparam ram_block1a24.port_b_data_out_clear = "none";
defparam ram_block1a24.port_b_data_out_clock = "none";
defparam ram_block1a24.port_b_data_width = 1;
defparam ram_block1a24.port_b_first_address = 0;
defparam ram_block1a24.port_b_first_bit_number = 24;
defparam ram_block1a24.port_b_last_address = 31;
defparam ram_block1a24.port_b_logical_ram_depth = 32;
defparam ram_block1a24.port_b_logical_ram_width = 32;
defparam ram_block1a24.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a24.port_b_read_enable_clock = "clock0";
defparam ram_block1a24.ram_block_type = "auto";

cyclonev_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_register_bank_a_module:first_nios2_system_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_voi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "old";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 5;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 31;
defparam ram_block1a0.port_a_logical_ram_depth = 32;
defparam ram_block1a0.port_a_logical_ram_width = 32;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock0";
defparam ram_block1a0.port_b_address_width = 5;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "none";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 31;
defparam ram_block1a0.port_b_logical_ram_depth = 32;
defparam ram_block1a0.port_b_logical_ram_width = 32;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock0";
defparam ram_block1a0.ram_block_type = "auto";

cyclonev_ram_block ram_block1a25(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[25]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a25_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a25.data_interleave_offset_in_bits = 1;
defparam ram_block1a25.data_interleave_width_in_bits = 1;
defparam ram_block1a25.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_register_bank_a_module:first_nios2_system_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_voi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a25.mixed_port_feed_through_mode = "old";
defparam ram_block1a25.operation_mode = "dual_port";
defparam ram_block1a25.port_a_address_clear = "none";
defparam ram_block1a25.port_a_address_width = 5;
defparam ram_block1a25.port_a_data_out_clear = "none";
defparam ram_block1a25.port_a_data_out_clock = "none";
defparam ram_block1a25.port_a_data_width = 1;
defparam ram_block1a25.port_a_first_address = 0;
defparam ram_block1a25.port_a_first_bit_number = 25;
defparam ram_block1a25.port_a_last_address = 31;
defparam ram_block1a25.port_a_logical_ram_depth = 32;
defparam ram_block1a25.port_a_logical_ram_width = 32;
defparam ram_block1a25.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a25.port_b_address_clear = "none";
defparam ram_block1a25.port_b_address_clock = "clock0";
defparam ram_block1a25.port_b_address_width = 5;
defparam ram_block1a25.port_b_data_out_clear = "none";
defparam ram_block1a25.port_b_data_out_clock = "none";
defparam ram_block1a25.port_b_data_width = 1;
defparam ram_block1a25.port_b_first_address = 0;
defparam ram_block1a25.port_b_first_bit_number = 25;
defparam ram_block1a25.port_b_last_address = 31;
defparam ram_block1a25.port_b_logical_ram_depth = 32;
defparam ram_block1a25.port_b_logical_ram_width = 32;
defparam ram_block1a25.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a25.port_b_read_enable_clock = "clock0";
defparam ram_block1a25.ram_block_type = "auto";

cyclonev_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_register_bank_a_module:first_nios2_system_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_voi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "old";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 5;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 31;
defparam ram_block1a2.port_a_logical_ram_depth = 32;
defparam ram_block1a2.port_a_logical_ram_width = 32;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock0";
defparam ram_block1a2.port_b_address_width = 5;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "none";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 31;
defparam ram_block1a2.port_b_logical_ram_depth = 32;
defparam ram_block1a2.port_b_logical_ram_width = 32;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock0";
defparam ram_block1a2.ram_block_type = "auto";

cyclonev_ram_block ram_block1a31(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a31_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a31.data_interleave_offset_in_bits = 1;
defparam ram_block1a31.data_interleave_width_in_bits = 1;
defparam ram_block1a31.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_register_bank_a_module:first_nios2_system_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_voi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a31.mixed_port_feed_through_mode = "old";
defparam ram_block1a31.operation_mode = "dual_port";
defparam ram_block1a31.port_a_address_clear = "none";
defparam ram_block1a31.port_a_address_width = 5;
defparam ram_block1a31.port_a_data_out_clear = "none";
defparam ram_block1a31.port_a_data_out_clock = "none";
defparam ram_block1a31.port_a_data_width = 1;
defparam ram_block1a31.port_a_first_address = 0;
defparam ram_block1a31.port_a_first_bit_number = 31;
defparam ram_block1a31.port_a_last_address = 31;
defparam ram_block1a31.port_a_logical_ram_depth = 32;
defparam ram_block1a31.port_a_logical_ram_width = 32;
defparam ram_block1a31.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a31.port_b_address_clear = "none";
defparam ram_block1a31.port_b_address_clock = "clock0";
defparam ram_block1a31.port_b_address_width = 5;
defparam ram_block1a31.port_b_data_out_clear = "none";
defparam ram_block1a31.port_b_data_out_clock = "none";
defparam ram_block1a31.port_b_data_width = 1;
defparam ram_block1a31.port_b_first_address = 0;
defparam ram_block1a31.port_b_first_bit_number = 31;
defparam ram_block1a31.port_b_last_address = 31;
defparam ram_block1a31.port_b_logical_ram_depth = 32;
defparam ram_block1a31.port_b_logical_ram_width = 32;
defparam ram_block1a31.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a31.port_b_read_enable_clock = "clock0";
defparam ram_block1a31.ram_block_type = "auto";

cyclonev_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_register_bank_a_module:first_nios2_system_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_voi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "old";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 5;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 31;
defparam ram_block1a7.port_a_logical_ram_depth = 32;
defparam ram_block1a7.port_a_logical_ram_width = 32;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock0";
defparam ram_block1a7.port_b_address_width = 5;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "none";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 31;
defparam ram_block1a7.port_b_logical_ram_depth = 32;
defparam ram_block1a7.port_b_logical_ram_width = 32;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock0";
defparam ram_block1a7.ram_block_type = "auto";

cyclonev_ram_block ram_block1a21(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a21_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_register_bank_a_module:first_nios2_system_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_voi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a21.mixed_port_feed_through_mode = "old";
defparam ram_block1a21.operation_mode = "dual_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 5;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 31;
defparam ram_block1a21.port_a_logical_ram_depth = 32;
defparam ram_block1a21.port_a_logical_ram_width = 32;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a21.port_b_address_clear = "none";
defparam ram_block1a21.port_b_address_clock = "clock0";
defparam ram_block1a21.port_b_address_width = 5;
defparam ram_block1a21.port_b_data_out_clear = "none";
defparam ram_block1a21.port_b_data_out_clock = "none";
defparam ram_block1a21.port_b_data_width = 1;
defparam ram_block1a21.port_b_first_address = 0;
defparam ram_block1a21.port_b_first_bit_number = 21;
defparam ram_block1a21.port_b_last_address = 31;
defparam ram_block1a21.port_b_logical_ram_depth = 32;
defparam ram_block1a21.port_b_logical_ram_width = 32;
defparam ram_block1a21.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a21.port_b_read_enable_clock = "clock0";
defparam ram_block1a21.ram_block_type = "auto";

cyclonev_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_register_bank_a_module:first_nios2_system_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_voi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "old";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 5;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 31;
defparam ram_block1a11.port_a_logical_ram_depth = 32;
defparam ram_block1a11.port_a_logical_ram_width = 32;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock0";
defparam ram_block1a11.port_b_address_width = 5;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "none";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 31;
defparam ram_block1a11.port_b_logical_ram_depth = 32;
defparam ram_block1a11.port_b_logical_ram_width = 32;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock0";
defparam ram_block1a11.ram_block_type = "auto";

cyclonev_ram_block ram_block1a28(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[28]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a28_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a28.data_interleave_offset_in_bits = 1;
defparam ram_block1a28.data_interleave_width_in_bits = 1;
defparam ram_block1a28.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_register_bank_a_module:first_nios2_system_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_voi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a28.mixed_port_feed_through_mode = "old";
defparam ram_block1a28.operation_mode = "dual_port";
defparam ram_block1a28.port_a_address_clear = "none";
defparam ram_block1a28.port_a_address_width = 5;
defparam ram_block1a28.port_a_data_out_clear = "none";
defparam ram_block1a28.port_a_data_out_clock = "none";
defparam ram_block1a28.port_a_data_width = 1;
defparam ram_block1a28.port_a_first_address = 0;
defparam ram_block1a28.port_a_first_bit_number = 28;
defparam ram_block1a28.port_a_last_address = 31;
defparam ram_block1a28.port_a_logical_ram_depth = 32;
defparam ram_block1a28.port_a_logical_ram_width = 32;
defparam ram_block1a28.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a28.port_b_address_clear = "none";
defparam ram_block1a28.port_b_address_clock = "clock0";
defparam ram_block1a28.port_b_address_width = 5;
defparam ram_block1a28.port_b_data_out_clear = "none";
defparam ram_block1a28.port_b_data_out_clock = "none";
defparam ram_block1a28.port_b_data_width = 1;
defparam ram_block1a28.port_b_first_address = 0;
defparam ram_block1a28.port_b_first_bit_number = 28;
defparam ram_block1a28.port_b_last_address = 31;
defparam ram_block1a28.port_b_logical_ram_depth = 32;
defparam ram_block1a28.port_b_logical_ram_width = 32;
defparam ram_block1a28.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a28.port_b_read_enable_clock = "clock0";
defparam ram_block1a28.ram_block_type = "auto";

cyclonev_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_register_bank_a_module:first_nios2_system_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_voi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "old";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 5;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 31;
defparam ram_block1a10.port_a_logical_ram_depth = 32;
defparam ram_block1a10.port_a_logical_ram_width = 32;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock0";
defparam ram_block1a10.port_b_address_width = 5;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "none";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 31;
defparam ram_block1a10.port_b_logical_ram_depth = 32;
defparam ram_block1a10.port_b_logical_ram_width = 32;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock0";
defparam ram_block1a10.ram_block_type = "auto";

cyclonev_ram_block ram_block1a27(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[27]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a27_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a27.data_interleave_offset_in_bits = 1;
defparam ram_block1a27.data_interleave_width_in_bits = 1;
defparam ram_block1a27.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_register_bank_a_module:first_nios2_system_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_voi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a27.mixed_port_feed_through_mode = "old";
defparam ram_block1a27.operation_mode = "dual_port";
defparam ram_block1a27.port_a_address_clear = "none";
defparam ram_block1a27.port_a_address_width = 5;
defparam ram_block1a27.port_a_data_out_clear = "none";
defparam ram_block1a27.port_a_data_out_clock = "none";
defparam ram_block1a27.port_a_data_width = 1;
defparam ram_block1a27.port_a_first_address = 0;
defparam ram_block1a27.port_a_first_bit_number = 27;
defparam ram_block1a27.port_a_last_address = 31;
defparam ram_block1a27.port_a_logical_ram_depth = 32;
defparam ram_block1a27.port_a_logical_ram_width = 32;
defparam ram_block1a27.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a27.port_b_address_clear = "none";
defparam ram_block1a27.port_b_address_clock = "clock0";
defparam ram_block1a27.port_b_address_width = 5;
defparam ram_block1a27.port_b_data_out_clear = "none";
defparam ram_block1a27.port_b_data_out_clock = "none";
defparam ram_block1a27.port_b_data_width = 1;
defparam ram_block1a27.port_b_first_address = 0;
defparam ram_block1a27.port_b_first_bit_number = 27;
defparam ram_block1a27.port_b_last_address = 31;
defparam ram_block1a27.port_b_logical_ram_depth = 32;
defparam ram_block1a27.port_b_logical_ram_width = 32;
defparam ram_block1a27.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a27.port_b_read_enable_clock = "clock0";
defparam ram_block1a27.ram_block_type = "auto";

cyclonev_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_register_bank_a_module:first_nios2_system_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_voi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "old";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 5;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 31;
defparam ram_block1a8.port_a_logical_ram_depth = 32;
defparam ram_block1a8.port_a_logical_ram_width = 32;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock0";
defparam ram_block1a8.port_b_address_width = 5;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "none";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 31;
defparam ram_block1a8.port_b_logical_ram_depth = 32;
defparam ram_block1a8.port_b_logical_ram_width = 32;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock0";
defparam ram_block1a8.ram_block_type = "auto";

cyclonev_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_register_bank_a_module:first_nios2_system_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_voi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "old";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 5;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 31;
defparam ram_block1a9.port_a_logical_ram_depth = 32;
defparam ram_block1a9.port_a_logical_ram_width = 32;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock0";
defparam ram_block1a9.port_b_address_width = 5;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "none";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 31;
defparam ram_block1a9.port_b_logical_ram_depth = 32;
defparam ram_block1a9.port_b_logical_ram_width = 32;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock0";
defparam ram_block1a9.ram_block_type = "auto";

cyclonev_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_register_bank_a_module:first_nios2_system_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_voi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "old";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 5;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 31;
defparam ram_block1a4.port_a_logical_ram_depth = 32;
defparam ram_block1a4.port_a_logical_ram_width = 32;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock0";
defparam ram_block1a4.port_b_address_width = 5;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "none";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 31;
defparam ram_block1a4.port_b_logical_ram_depth = 32;
defparam ram_block1a4.port_b_logical_ram_width = 32;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock0";
defparam ram_block1a4.ram_block_type = "auto";

cyclonev_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_register_bank_a_module:first_nios2_system_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_voi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "old";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 5;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 31;
defparam ram_block1a5.port_a_logical_ram_depth = 32;
defparam ram_block1a5.port_a_logical_ram_width = 32;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock0";
defparam ram_block1a5.port_b_address_width = 5;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "none";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 31;
defparam ram_block1a5.port_b_logical_ram_depth = 32;
defparam ram_block1a5.port_b_logical_ram_width = 32;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock0";
defparam ram_block1a5.ram_block_type = "auto";

cyclonev_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_register_bank_a_module:first_nios2_system_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_voi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "old";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 5;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 31;
defparam ram_block1a6.port_a_logical_ram_depth = 32;
defparam ram_block1a6.port_a_logical_ram_width = 32;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock0";
defparam ram_block1a6.port_b_address_width = 5;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "none";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 31;
defparam ram_block1a6.port_b_logical_ram_depth = 32;
defparam ram_block1a6.port_b_logical_ram_width = 32;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock0";
defparam ram_block1a6.ram_block_type = "auto";

cyclonev_ram_block ram_block1a26(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[26]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a26_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a26.data_interleave_offset_in_bits = 1;
defparam ram_block1a26.data_interleave_width_in_bits = 1;
defparam ram_block1a26.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_register_bank_a_module:first_nios2_system_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_voi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a26.mixed_port_feed_through_mode = "old";
defparam ram_block1a26.operation_mode = "dual_port";
defparam ram_block1a26.port_a_address_clear = "none";
defparam ram_block1a26.port_a_address_width = 5;
defparam ram_block1a26.port_a_data_out_clear = "none";
defparam ram_block1a26.port_a_data_out_clock = "none";
defparam ram_block1a26.port_a_data_width = 1;
defparam ram_block1a26.port_a_first_address = 0;
defparam ram_block1a26.port_a_first_bit_number = 26;
defparam ram_block1a26.port_a_last_address = 31;
defparam ram_block1a26.port_a_logical_ram_depth = 32;
defparam ram_block1a26.port_a_logical_ram_width = 32;
defparam ram_block1a26.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a26.port_b_address_clear = "none";
defparam ram_block1a26.port_b_address_clock = "clock0";
defparam ram_block1a26.port_b_address_width = 5;
defparam ram_block1a26.port_b_data_out_clear = "none";
defparam ram_block1a26.port_b_data_out_clock = "none";
defparam ram_block1a26.port_b_data_width = 1;
defparam ram_block1a26.port_b_first_address = 0;
defparam ram_block1a26.port_b_first_bit_number = 26;
defparam ram_block1a26.port_b_last_address = 31;
defparam ram_block1a26.port_b_logical_ram_depth = 32;
defparam ram_block1a26.port_b_logical_ram_width = 32;
defparam ram_block1a26.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a26.port_b_read_enable_clock = "clock0";
defparam ram_block1a26.ram_block_type = "auto";

cyclonev_ram_block ram_block1a20(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a20_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_register_bank_a_module:first_nios2_system_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_voi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a20.mixed_port_feed_through_mode = "old";
defparam ram_block1a20.operation_mode = "dual_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 5;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 31;
defparam ram_block1a20.port_a_logical_ram_depth = 32;
defparam ram_block1a20.port_a_logical_ram_width = 32;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a20.port_b_address_clear = "none";
defparam ram_block1a20.port_b_address_clock = "clock0";
defparam ram_block1a20.port_b_address_width = 5;
defparam ram_block1a20.port_b_data_out_clear = "none";
defparam ram_block1a20.port_b_data_out_clock = "none";
defparam ram_block1a20.port_b_data_width = 1;
defparam ram_block1a20.port_b_first_address = 0;
defparam ram_block1a20.port_b_first_bit_number = 20;
defparam ram_block1a20.port_b_last_address = 31;
defparam ram_block1a20.port_b_logical_ram_depth = 32;
defparam ram_block1a20.port_b_logical_ram_width = 32;
defparam ram_block1a20.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a20.port_b_read_enable_clock = "clock0";
defparam ram_block1a20.ram_block_type = "auto";

cyclonev_ram_block ram_block1a19(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a19_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_register_bank_a_module:first_nios2_system_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_voi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a19.mixed_port_feed_through_mode = "old";
defparam ram_block1a19.operation_mode = "dual_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 5;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 31;
defparam ram_block1a19.port_a_logical_ram_depth = 32;
defparam ram_block1a19.port_a_logical_ram_width = 32;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a19.port_b_address_clear = "none";
defparam ram_block1a19.port_b_address_clock = "clock0";
defparam ram_block1a19.port_b_address_width = 5;
defparam ram_block1a19.port_b_data_out_clear = "none";
defparam ram_block1a19.port_b_data_out_clock = "none";
defparam ram_block1a19.port_b_data_width = 1;
defparam ram_block1a19.port_b_first_address = 0;
defparam ram_block1a19.port_b_first_bit_number = 19;
defparam ram_block1a19.port_b_last_address = 31;
defparam ram_block1a19.port_b_logical_ram_depth = 32;
defparam ram_block1a19.port_b_logical_ram_width = 32;
defparam ram_block1a19.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a19.port_b_read_enable_clock = "clock0";
defparam ram_block1a19.ram_block_type = "auto";

cyclonev_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_register_bank_a_module:first_nios2_system_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_voi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "old";
defparam ram_block1a17.operation_mode = "dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 5;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 31;
defparam ram_block1a17.port_a_logical_ram_depth = 32;
defparam ram_block1a17.port_a_logical_ram_width = 32;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a17.port_b_address_clear = "none";
defparam ram_block1a17.port_b_address_clock = "clock0";
defparam ram_block1a17.port_b_address_width = 5;
defparam ram_block1a17.port_b_data_out_clear = "none";
defparam ram_block1a17.port_b_data_out_clock = "none";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 31;
defparam ram_block1a17.port_b_logical_ram_depth = 32;
defparam ram_block1a17.port_b_logical_ram_width = 32;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock0";
defparam ram_block1a17.ram_block_type = "auto";

cyclonev_ram_block ram_block1a30(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[30]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a30_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a30.data_interleave_offset_in_bits = 1;
defparam ram_block1a30.data_interleave_width_in_bits = 1;
defparam ram_block1a30.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_register_bank_a_module:first_nios2_system_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_voi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a30.mixed_port_feed_through_mode = "old";
defparam ram_block1a30.operation_mode = "dual_port";
defparam ram_block1a30.port_a_address_clear = "none";
defparam ram_block1a30.port_a_address_width = 5;
defparam ram_block1a30.port_a_data_out_clear = "none";
defparam ram_block1a30.port_a_data_out_clock = "none";
defparam ram_block1a30.port_a_data_width = 1;
defparam ram_block1a30.port_a_first_address = 0;
defparam ram_block1a30.port_a_first_bit_number = 30;
defparam ram_block1a30.port_a_last_address = 31;
defparam ram_block1a30.port_a_logical_ram_depth = 32;
defparam ram_block1a30.port_a_logical_ram_width = 32;
defparam ram_block1a30.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a30.port_b_address_clear = "none";
defparam ram_block1a30.port_b_address_clock = "clock0";
defparam ram_block1a30.port_b_address_width = 5;
defparam ram_block1a30.port_b_data_out_clear = "none";
defparam ram_block1a30.port_b_data_out_clock = "none";
defparam ram_block1a30.port_b_data_width = 1;
defparam ram_block1a30.port_b_first_address = 0;
defparam ram_block1a30.port_b_first_bit_number = 30;
defparam ram_block1a30.port_b_last_address = 31;
defparam ram_block1a30.port_b_logical_ram_depth = 32;
defparam ram_block1a30.port_b_logical_ram_width = 32;
defparam ram_block1a30.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a30.port_b_read_enable_clock = "clock0";
defparam ram_block1a30.ram_block_type = "auto";

cyclonev_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_register_bank_a_module:first_nios2_system_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_voi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "old";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 5;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 31;
defparam ram_block1a1.port_a_logical_ram_depth = 32;
defparam ram_block1a1.port_a_logical_ram_width = 32;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock0";
defparam ram_block1a1.port_b_address_width = 5;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "none";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 31;
defparam ram_block1a1.port_b_logical_ram_depth = 32;
defparam ram_block1a1.port_b_logical_ram_width = 32;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock0";
defparam ram_block1a1.ram_block_type = "auto";

cyclonev_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_register_bank_a_module:first_nios2_system_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_voi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "old";
defparam ram_block1a18.operation_mode = "dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 5;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 31;
defparam ram_block1a18.port_a_logical_ram_depth = 32;
defparam ram_block1a18.port_a_logical_ram_width = 32;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a18.port_b_address_clear = "none";
defparam ram_block1a18.port_b_address_clock = "clock0";
defparam ram_block1a18.port_b_address_width = 5;
defparam ram_block1a18.port_b_data_out_clear = "none";
defparam ram_block1a18.port_b_data_out_clock = "none";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 31;
defparam ram_block1a18.port_b_logical_ram_depth = 32;
defparam ram_block1a18.port_b_logical_ram_width = 32;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock0";
defparam ram_block1a18.ram_block_type = "auto";

cyclonev_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_register_bank_a_module:first_nios2_system_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_voi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "old";
defparam ram_block1a16.operation_mode = "dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 5;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 31;
defparam ram_block1a16.port_a_logical_ram_depth = 32;
defparam ram_block1a16.port_a_logical_ram_width = 32;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a16.port_b_address_clear = "none";
defparam ram_block1a16.port_b_address_clock = "clock0";
defparam ram_block1a16.port_b_address_width = 5;
defparam ram_block1a16.port_b_data_out_clear = "none";
defparam ram_block1a16.port_b_data_out_clock = "none";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 31;
defparam ram_block1a16.port_b_logical_ram_depth = 32;
defparam ram_block1a16.port_b_logical_ram_width = 32;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock0";
defparam ram_block1a16.ram_block_type = "auto";

cyclonev_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_register_bank_a_module:first_nios2_system_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_voi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "old";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 5;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 31;
defparam ram_block1a15.port_a_logical_ram_depth = 32;
defparam ram_block1a15.port_a_logical_ram_width = 32;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock0";
defparam ram_block1a15.port_b_address_width = 5;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "none";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 31;
defparam ram_block1a15.port_b_logical_ram_depth = 32;
defparam ram_block1a15.port_b_logical_ram_width = 32;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock0";
defparam ram_block1a15.ram_block_type = "auto";

cyclonev_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_register_bank_a_module:first_nios2_system_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_voi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "old";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 5;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 31;
defparam ram_block1a12.port_a_logical_ram_depth = 32;
defparam ram_block1a12.port_a_logical_ram_width = 32;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock0";
defparam ram_block1a12.port_b_address_width = 5;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "none";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 31;
defparam ram_block1a12.port_b_logical_ram_depth = 32;
defparam ram_block1a12.port_b_logical_ram_width = 32;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock0";
defparam ram_block1a12.ram_block_type = "auto";

cyclonev_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_register_bank_a_module:first_nios2_system_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_voi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "old";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 5;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 31;
defparam ram_block1a13.port_a_logical_ram_depth = 32;
defparam ram_block1a13.port_a_logical_ram_width = 32;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock0";
defparam ram_block1a13.port_b_address_width = 5;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "none";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 31;
defparam ram_block1a13.port_b_logical_ram_depth = 32;
defparam ram_block1a13.port_b_logical_ram_width = 32;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock0";
defparam ram_block1a13.ram_block_type = "auto";

cyclonev_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_register_bank_a_module:first_nios2_system_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_voi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "old";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 5;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 31;
defparam ram_block1a14.port_a_logical_ram_depth = 32;
defparam ram_block1a14.port_a_logical_ram_width = 32;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock0";
defparam ram_block1a14.port_b_address_width = 5;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "none";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 31;
defparam ram_block1a14.port_b_logical_ram_depth = 32;
defparam ram_block1a14.port_b_logical_ram_width = 32;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock0";
defparam ram_block1a14.ram_block_type = "auto";

cyclonev_ram_block ram_block1a29(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[29]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a29_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a29.data_interleave_offset_in_bits = 1;
defparam ram_block1a29.data_interleave_width_in_bits = 1;
defparam ram_block1a29.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_register_bank_a_module:first_nios2_system_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_voi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a29.mixed_port_feed_through_mode = "old";
defparam ram_block1a29.operation_mode = "dual_port";
defparam ram_block1a29.port_a_address_clear = "none";
defparam ram_block1a29.port_a_address_width = 5;
defparam ram_block1a29.port_a_data_out_clear = "none";
defparam ram_block1a29.port_a_data_out_clock = "none";
defparam ram_block1a29.port_a_data_width = 1;
defparam ram_block1a29.port_a_first_address = 0;
defparam ram_block1a29.port_a_first_bit_number = 29;
defparam ram_block1a29.port_a_last_address = 31;
defparam ram_block1a29.port_a_logical_ram_depth = 32;
defparam ram_block1a29.port_a_logical_ram_width = 32;
defparam ram_block1a29.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a29.port_b_address_clear = "none";
defparam ram_block1a29.port_b_address_clock = "clock0";
defparam ram_block1a29.port_b_address_width = 5;
defparam ram_block1a29.port_b_data_out_clear = "none";
defparam ram_block1a29.port_b_data_out_clock = "none";
defparam ram_block1a29.port_b_data_width = 1;
defparam ram_block1a29.port_b_first_address = 0;
defparam ram_block1a29.port_b_first_bit_number = 29;
defparam ram_block1a29.port_b_last_address = 31;
defparam ram_block1a29.port_b_logical_ram_depth = 32;
defparam ram_block1a29.port_b_logical_ram_width = 32;
defparam ram_block1a29.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a29.port_b_read_enable_clock = "clock0";
defparam ram_block1a29.ram_block_type = "auto";

endmodule

module first_nios2_system_first_nios2_system_cpu_cpu_register_bank_b_module (
	q_b_0,
	q_b_1,
	q_b_2,
	q_b_3,
	q_b_4,
	q_b_5,
	q_b_6,
	q_b_7,
	q_b_22,
	q_b_23,
	q_b_24,
	q_b_25,
	q_b_31,
	q_b_21,
	q_b_11,
	q_b_28,
	q_b_10,
	q_b_27,
	q_b_8,
	q_b_9,
	q_b_26,
	q_b_20,
	q_b_19,
	q_b_17,
	q_b_30,
	q_b_18,
	q_b_16,
	q_b_15,
	q_b_12,
	q_b_13,
	q_b_14,
	q_b_29,
	A_wr_data_unfiltered_0,
	A_wr_data_unfiltered_1,
	A_wr_data_unfiltered_2,
	A_wr_data_unfiltered_3,
	A_wr_data_unfiltered_4,
	A_wr_data_unfiltered_5,
	A_wr_data_unfiltered_6,
	A_wr_data_unfiltered_7,
	A_wr_data_unfiltered_22,
	A_wr_data_unfiltered_23,
	A_wr_data_unfiltered_24,
	A_wr_data_unfiltered_25,
	A_wr_data_unfiltered_31,
	A_wr_data_unfiltered_21,
	A_wr_data_unfiltered_11,
	A_wr_data_unfiltered_28,
	A_wr_data_unfiltered_10,
	A_wr_data_unfiltered_27,
	A_wr_data_unfiltered_8,
	A_wr_data_unfiltered_9,
	A_wr_data_unfiltered_26,
	A_wr_data_unfiltered_20,
	A_wr_data_unfiltered_19,
	A_wr_data_unfiltered_17,
	A_wr_data_unfiltered_30,
	A_wr_data_unfiltered_18,
	A_wr_data_unfiltered_16,
	A_wr_data_unfiltered_15,
	A_wr_data_unfiltered_12,
	A_wr_data_unfiltered_13,
	A_wr_data_unfiltered_14,
	A_wr_data_unfiltered_29,
	A_wr_dst_reg,
	A_dst_regnum,
	A_dst_regnum1,
	A_dst_regnum2,
	A_dst_regnum3,
	A_dst_regnum4,
	rf_b_rd_port_addr_0,
	rf_b_rd_port_addr_1,
	rf_b_rd_port_addr_2,
	rf_b_rd_port_addr_3,
	rf_b_rd_port_addr_4,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_0;
output 	q_b_1;
output 	q_b_2;
output 	q_b_3;
output 	q_b_4;
output 	q_b_5;
output 	q_b_6;
output 	q_b_7;
output 	q_b_22;
output 	q_b_23;
output 	q_b_24;
output 	q_b_25;
output 	q_b_31;
output 	q_b_21;
output 	q_b_11;
output 	q_b_28;
output 	q_b_10;
output 	q_b_27;
output 	q_b_8;
output 	q_b_9;
output 	q_b_26;
output 	q_b_20;
output 	q_b_19;
output 	q_b_17;
output 	q_b_30;
output 	q_b_18;
output 	q_b_16;
output 	q_b_15;
output 	q_b_12;
output 	q_b_13;
output 	q_b_14;
output 	q_b_29;
input 	A_wr_data_unfiltered_0;
input 	A_wr_data_unfiltered_1;
input 	A_wr_data_unfiltered_2;
input 	A_wr_data_unfiltered_3;
input 	A_wr_data_unfiltered_4;
input 	A_wr_data_unfiltered_5;
input 	A_wr_data_unfiltered_6;
input 	A_wr_data_unfiltered_7;
input 	A_wr_data_unfiltered_22;
input 	A_wr_data_unfiltered_23;
input 	A_wr_data_unfiltered_24;
input 	A_wr_data_unfiltered_25;
input 	A_wr_data_unfiltered_31;
input 	A_wr_data_unfiltered_21;
input 	A_wr_data_unfiltered_11;
input 	A_wr_data_unfiltered_28;
input 	A_wr_data_unfiltered_10;
input 	A_wr_data_unfiltered_27;
input 	A_wr_data_unfiltered_8;
input 	A_wr_data_unfiltered_9;
input 	A_wr_data_unfiltered_26;
input 	A_wr_data_unfiltered_20;
input 	A_wr_data_unfiltered_19;
input 	A_wr_data_unfiltered_17;
input 	A_wr_data_unfiltered_30;
input 	A_wr_data_unfiltered_18;
input 	A_wr_data_unfiltered_16;
input 	A_wr_data_unfiltered_15;
input 	A_wr_data_unfiltered_12;
input 	A_wr_data_unfiltered_13;
input 	A_wr_data_unfiltered_14;
input 	A_wr_data_unfiltered_29;
input 	A_wr_dst_reg;
input 	A_dst_regnum;
input 	A_dst_regnum1;
input 	A_dst_regnum2;
input 	A_dst_regnum3;
input 	A_dst_regnum4;
input 	rf_b_rd_port_addr_0;
input 	rf_b_rd_port_addr_1;
input 	rf_b_rd_port_addr_2;
input 	rf_b_rd_port_addr_3;
input 	rf_b_rd_port_addr_4;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



first_nios2_system_altsyncram_6 the_altsyncram(
	.q_b({q_b_31,q_b_30,q_b_29,q_b_28,q_b_27,q_b_26,q_b_25,q_b_24,q_b_23,q_b_22,q_b_21,q_b_20,q_b_19,q_b_18,q_b_17,q_b_16,q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.data_a({A_wr_data_unfiltered_31,A_wr_data_unfiltered_30,A_wr_data_unfiltered_29,A_wr_data_unfiltered_28,A_wr_data_unfiltered_27,A_wr_data_unfiltered_26,A_wr_data_unfiltered_25,A_wr_data_unfiltered_24,A_wr_data_unfiltered_23,A_wr_data_unfiltered_22,A_wr_data_unfiltered_21,
A_wr_data_unfiltered_20,A_wr_data_unfiltered_19,A_wr_data_unfiltered_18,A_wr_data_unfiltered_17,A_wr_data_unfiltered_16,A_wr_data_unfiltered_15,A_wr_data_unfiltered_14,A_wr_data_unfiltered_13,A_wr_data_unfiltered_12,A_wr_data_unfiltered_11,A_wr_data_unfiltered_10,
A_wr_data_unfiltered_9,A_wr_data_unfiltered_8,A_wr_data_unfiltered_7,A_wr_data_unfiltered_6,A_wr_data_unfiltered_5,A_wr_data_unfiltered_4,A_wr_data_unfiltered_3,A_wr_data_unfiltered_2,A_wr_data_unfiltered_1,A_wr_data_unfiltered_0}),
	.wren_a(A_wr_dst_reg),
	.address_a({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,A_dst_regnum4,A_dst_regnum3,A_dst_regnum2,A_dst_regnum1,A_dst_regnum}),
	.address_b({gnd,gnd,gnd,gnd,rf_b_rd_port_addr_4,rf_b_rd_port_addr_3,rf_b_rd_port_addr_2,rf_b_rd_port_addr_1,rf_b_rd_port_addr_0}),
	.clock0(clk_clk));

endmodule

module first_nios2_system_altsyncram_6 (
	q_b,
	data_a,
	wren_a,
	address_a,
	address_b,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_b;
input 	[31:0] data_a;
input 	wren_a;
input 	[12:0] address_a;
input 	[8:0] address_b;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



first_nios2_system_altsyncram_voi1_1 auto_generated(
	.q_b({q_b[31],q_b[30],q_b[29],q_b[28],q_b[27],q_b[26],q_b[25],q_b[24],q_b[23],q_b[22],q_b[21],q_b[20],q_b[19],q_b[18],q_b[17],q_b[16],q_b[15],q_b[14],q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.data_a({data_a[31],data_a[30],data_a[29],data_a[28],data_a[27],data_a[26],data_a[25],data_a[24],data_a[23],data_a[22],data_a[21],data_a[20],data_a[19],data_a[18],data_a[17],data_a[16],data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.wren_a(wren_a),
	.address_a({address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.address_b({address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.clock0(clock0));

endmodule

module first_nios2_system_altsyncram_voi1_1 (
	q_b,
	data_a,
	wren_a,
	address_a,
	address_b,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_b;
input 	[31:0] data_a;
input 	wren_a;
input 	[4:0] address_a;
input 	[4:0] address_b;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a22_PORTBDATAOUT_bus;
wire [143:0] ram_block1a23_PORTBDATAOUT_bus;
wire [143:0] ram_block1a24_PORTBDATAOUT_bus;
wire [143:0] ram_block1a25_PORTBDATAOUT_bus;
wire [143:0] ram_block1a31_PORTBDATAOUT_bus;
wire [143:0] ram_block1a21_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a28_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a27_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a26_PORTBDATAOUT_bus;
wire [143:0] ram_block1a20_PORTBDATAOUT_bus;
wire [143:0] ram_block1a19_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;
wire [143:0] ram_block1a30_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a29_PORTBDATAOUT_bus;

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[22] = ram_block1a22_PORTBDATAOUT_bus[0];

assign q_b[23] = ram_block1a23_PORTBDATAOUT_bus[0];

assign q_b[24] = ram_block1a24_PORTBDATAOUT_bus[0];

assign q_b[25] = ram_block1a25_PORTBDATAOUT_bus[0];

assign q_b[31] = ram_block1a31_PORTBDATAOUT_bus[0];

assign q_b[21] = ram_block1a21_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[28] = ram_block1a28_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[27] = ram_block1a27_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[26] = ram_block1a26_PORTBDATAOUT_bus[0];

assign q_b[20] = ram_block1a20_PORTBDATAOUT_bus[0];

assign q_b[19] = ram_block1a19_PORTBDATAOUT_bus[0];

assign q_b[17] = ram_block1a17_PORTBDATAOUT_bus[0];

assign q_b[30] = ram_block1a30_PORTBDATAOUT_bus[0];

assign q_b[18] = ram_block1a18_PORTBDATAOUT_bus[0];

assign q_b[16] = ram_block1a16_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[29] = ram_block1a29_PORTBDATAOUT_bus[0];

cyclonev_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_register_bank_b_module:first_nios2_system_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_voi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "old";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 5;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 31;
defparam ram_block1a0.port_a_logical_ram_depth = 32;
defparam ram_block1a0.port_a_logical_ram_width = 32;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock0";
defparam ram_block1a0.port_b_address_width = 5;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "none";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 31;
defparam ram_block1a0.port_b_logical_ram_depth = 32;
defparam ram_block1a0.port_b_logical_ram_width = 32;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock0";
defparam ram_block1a0.ram_block_type = "auto";

cyclonev_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_register_bank_b_module:first_nios2_system_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_voi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "old";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 5;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 31;
defparam ram_block1a1.port_a_logical_ram_depth = 32;
defparam ram_block1a1.port_a_logical_ram_width = 32;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock0";
defparam ram_block1a1.port_b_address_width = 5;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "none";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 31;
defparam ram_block1a1.port_b_logical_ram_depth = 32;
defparam ram_block1a1.port_b_logical_ram_width = 32;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock0";
defparam ram_block1a1.ram_block_type = "auto";

cyclonev_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_register_bank_b_module:first_nios2_system_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_voi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "old";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 5;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 31;
defparam ram_block1a2.port_a_logical_ram_depth = 32;
defparam ram_block1a2.port_a_logical_ram_width = 32;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock0";
defparam ram_block1a2.port_b_address_width = 5;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "none";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 31;
defparam ram_block1a2.port_b_logical_ram_depth = 32;
defparam ram_block1a2.port_b_logical_ram_width = 32;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock0";
defparam ram_block1a2.ram_block_type = "auto";

cyclonev_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_register_bank_b_module:first_nios2_system_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_voi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "old";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 5;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 31;
defparam ram_block1a3.port_a_logical_ram_depth = 32;
defparam ram_block1a3.port_a_logical_ram_width = 32;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock0";
defparam ram_block1a3.port_b_address_width = 5;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "none";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 31;
defparam ram_block1a3.port_b_logical_ram_depth = 32;
defparam ram_block1a3.port_b_logical_ram_width = 32;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock0";
defparam ram_block1a3.ram_block_type = "auto";

cyclonev_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_register_bank_b_module:first_nios2_system_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_voi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "old";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 5;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 31;
defparam ram_block1a4.port_a_logical_ram_depth = 32;
defparam ram_block1a4.port_a_logical_ram_width = 32;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock0";
defparam ram_block1a4.port_b_address_width = 5;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "none";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 31;
defparam ram_block1a4.port_b_logical_ram_depth = 32;
defparam ram_block1a4.port_b_logical_ram_width = 32;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock0";
defparam ram_block1a4.ram_block_type = "auto";

cyclonev_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_register_bank_b_module:first_nios2_system_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_voi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "old";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 5;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 31;
defparam ram_block1a5.port_a_logical_ram_depth = 32;
defparam ram_block1a5.port_a_logical_ram_width = 32;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock0";
defparam ram_block1a5.port_b_address_width = 5;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "none";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 31;
defparam ram_block1a5.port_b_logical_ram_depth = 32;
defparam ram_block1a5.port_b_logical_ram_width = 32;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock0";
defparam ram_block1a5.ram_block_type = "auto";

cyclonev_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_register_bank_b_module:first_nios2_system_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_voi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "old";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 5;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 31;
defparam ram_block1a6.port_a_logical_ram_depth = 32;
defparam ram_block1a6.port_a_logical_ram_width = 32;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock0";
defparam ram_block1a6.port_b_address_width = 5;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "none";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 31;
defparam ram_block1a6.port_b_logical_ram_depth = 32;
defparam ram_block1a6.port_b_logical_ram_width = 32;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock0";
defparam ram_block1a6.ram_block_type = "auto";

cyclonev_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_register_bank_b_module:first_nios2_system_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_voi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "old";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 5;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 31;
defparam ram_block1a7.port_a_logical_ram_depth = 32;
defparam ram_block1a7.port_a_logical_ram_width = 32;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock0";
defparam ram_block1a7.port_b_address_width = 5;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "none";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 31;
defparam ram_block1a7.port_b_logical_ram_depth = 32;
defparam ram_block1a7.port_b_logical_ram_width = 32;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock0";
defparam ram_block1a7.ram_block_type = "auto";

cyclonev_ram_block ram_block1a22(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[22]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a22_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a22.data_interleave_offset_in_bits = 1;
defparam ram_block1a22.data_interleave_width_in_bits = 1;
defparam ram_block1a22.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_register_bank_b_module:first_nios2_system_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_voi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a22.mixed_port_feed_through_mode = "old";
defparam ram_block1a22.operation_mode = "dual_port";
defparam ram_block1a22.port_a_address_clear = "none";
defparam ram_block1a22.port_a_address_width = 5;
defparam ram_block1a22.port_a_data_out_clear = "none";
defparam ram_block1a22.port_a_data_out_clock = "none";
defparam ram_block1a22.port_a_data_width = 1;
defparam ram_block1a22.port_a_first_address = 0;
defparam ram_block1a22.port_a_first_bit_number = 22;
defparam ram_block1a22.port_a_last_address = 31;
defparam ram_block1a22.port_a_logical_ram_depth = 32;
defparam ram_block1a22.port_a_logical_ram_width = 32;
defparam ram_block1a22.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a22.port_b_address_clear = "none";
defparam ram_block1a22.port_b_address_clock = "clock0";
defparam ram_block1a22.port_b_address_width = 5;
defparam ram_block1a22.port_b_data_out_clear = "none";
defparam ram_block1a22.port_b_data_out_clock = "none";
defparam ram_block1a22.port_b_data_width = 1;
defparam ram_block1a22.port_b_first_address = 0;
defparam ram_block1a22.port_b_first_bit_number = 22;
defparam ram_block1a22.port_b_last_address = 31;
defparam ram_block1a22.port_b_logical_ram_depth = 32;
defparam ram_block1a22.port_b_logical_ram_width = 32;
defparam ram_block1a22.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a22.port_b_read_enable_clock = "clock0";
defparam ram_block1a22.ram_block_type = "auto";

cyclonev_ram_block ram_block1a23(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[23]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a23_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a23.data_interleave_offset_in_bits = 1;
defparam ram_block1a23.data_interleave_width_in_bits = 1;
defparam ram_block1a23.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_register_bank_b_module:first_nios2_system_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_voi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a23.mixed_port_feed_through_mode = "old";
defparam ram_block1a23.operation_mode = "dual_port";
defparam ram_block1a23.port_a_address_clear = "none";
defparam ram_block1a23.port_a_address_width = 5;
defparam ram_block1a23.port_a_data_out_clear = "none";
defparam ram_block1a23.port_a_data_out_clock = "none";
defparam ram_block1a23.port_a_data_width = 1;
defparam ram_block1a23.port_a_first_address = 0;
defparam ram_block1a23.port_a_first_bit_number = 23;
defparam ram_block1a23.port_a_last_address = 31;
defparam ram_block1a23.port_a_logical_ram_depth = 32;
defparam ram_block1a23.port_a_logical_ram_width = 32;
defparam ram_block1a23.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a23.port_b_address_clear = "none";
defparam ram_block1a23.port_b_address_clock = "clock0";
defparam ram_block1a23.port_b_address_width = 5;
defparam ram_block1a23.port_b_data_out_clear = "none";
defparam ram_block1a23.port_b_data_out_clock = "none";
defparam ram_block1a23.port_b_data_width = 1;
defparam ram_block1a23.port_b_first_address = 0;
defparam ram_block1a23.port_b_first_bit_number = 23;
defparam ram_block1a23.port_b_last_address = 31;
defparam ram_block1a23.port_b_logical_ram_depth = 32;
defparam ram_block1a23.port_b_logical_ram_width = 32;
defparam ram_block1a23.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a23.port_b_read_enable_clock = "clock0";
defparam ram_block1a23.ram_block_type = "auto";

cyclonev_ram_block ram_block1a24(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[24]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a24_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a24.data_interleave_offset_in_bits = 1;
defparam ram_block1a24.data_interleave_width_in_bits = 1;
defparam ram_block1a24.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_register_bank_b_module:first_nios2_system_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_voi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a24.mixed_port_feed_through_mode = "old";
defparam ram_block1a24.operation_mode = "dual_port";
defparam ram_block1a24.port_a_address_clear = "none";
defparam ram_block1a24.port_a_address_width = 5;
defparam ram_block1a24.port_a_data_out_clear = "none";
defparam ram_block1a24.port_a_data_out_clock = "none";
defparam ram_block1a24.port_a_data_width = 1;
defparam ram_block1a24.port_a_first_address = 0;
defparam ram_block1a24.port_a_first_bit_number = 24;
defparam ram_block1a24.port_a_last_address = 31;
defparam ram_block1a24.port_a_logical_ram_depth = 32;
defparam ram_block1a24.port_a_logical_ram_width = 32;
defparam ram_block1a24.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a24.port_b_address_clear = "none";
defparam ram_block1a24.port_b_address_clock = "clock0";
defparam ram_block1a24.port_b_address_width = 5;
defparam ram_block1a24.port_b_data_out_clear = "none";
defparam ram_block1a24.port_b_data_out_clock = "none";
defparam ram_block1a24.port_b_data_width = 1;
defparam ram_block1a24.port_b_first_address = 0;
defparam ram_block1a24.port_b_first_bit_number = 24;
defparam ram_block1a24.port_b_last_address = 31;
defparam ram_block1a24.port_b_logical_ram_depth = 32;
defparam ram_block1a24.port_b_logical_ram_width = 32;
defparam ram_block1a24.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a24.port_b_read_enable_clock = "clock0";
defparam ram_block1a24.ram_block_type = "auto";

cyclonev_ram_block ram_block1a25(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[25]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a25_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a25.data_interleave_offset_in_bits = 1;
defparam ram_block1a25.data_interleave_width_in_bits = 1;
defparam ram_block1a25.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_register_bank_b_module:first_nios2_system_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_voi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a25.mixed_port_feed_through_mode = "old";
defparam ram_block1a25.operation_mode = "dual_port";
defparam ram_block1a25.port_a_address_clear = "none";
defparam ram_block1a25.port_a_address_width = 5;
defparam ram_block1a25.port_a_data_out_clear = "none";
defparam ram_block1a25.port_a_data_out_clock = "none";
defparam ram_block1a25.port_a_data_width = 1;
defparam ram_block1a25.port_a_first_address = 0;
defparam ram_block1a25.port_a_first_bit_number = 25;
defparam ram_block1a25.port_a_last_address = 31;
defparam ram_block1a25.port_a_logical_ram_depth = 32;
defparam ram_block1a25.port_a_logical_ram_width = 32;
defparam ram_block1a25.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a25.port_b_address_clear = "none";
defparam ram_block1a25.port_b_address_clock = "clock0";
defparam ram_block1a25.port_b_address_width = 5;
defparam ram_block1a25.port_b_data_out_clear = "none";
defparam ram_block1a25.port_b_data_out_clock = "none";
defparam ram_block1a25.port_b_data_width = 1;
defparam ram_block1a25.port_b_first_address = 0;
defparam ram_block1a25.port_b_first_bit_number = 25;
defparam ram_block1a25.port_b_last_address = 31;
defparam ram_block1a25.port_b_logical_ram_depth = 32;
defparam ram_block1a25.port_b_logical_ram_width = 32;
defparam ram_block1a25.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a25.port_b_read_enable_clock = "clock0";
defparam ram_block1a25.ram_block_type = "auto";

cyclonev_ram_block ram_block1a31(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a31_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a31.data_interleave_offset_in_bits = 1;
defparam ram_block1a31.data_interleave_width_in_bits = 1;
defparam ram_block1a31.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_register_bank_b_module:first_nios2_system_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_voi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a31.mixed_port_feed_through_mode = "old";
defparam ram_block1a31.operation_mode = "dual_port";
defparam ram_block1a31.port_a_address_clear = "none";
defparam ram_block1a31.port_a_address_width = 5;
defparam ram_block1a31.port_a_data_out_clear = "none";
defparam ram_block1a31.port_a_data_out_clock = "none";
defparam ram_block1a31.port_a_data_width = 1;
defparam ram_block1a31.port_a_first_address = 0;
defparam ram_block1a31.port_a_first_bit_number = 31;
defparam ram_block1a31.port_a_last_address = 31;
defparam ram_block1a31.port_a_logical_ram_depth = 32;
defparam ram_block1a31.port_a_logical_ram_width = 32;
defparam ram_block1a31.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a31.port_b_address_clear = "none";
defparam ram_block1a31.port_b_address_clock = "clock0";
defparam ram_block1a31.port_b_address_width = 5;
defparam ram_block1a31.port_b_data_out_clear = "none";
defparam ram_block1a31.port_b_data_out_clock = "none";
defparam ram_block1a31.port_b_data_width = 1;
defparam ram_block1a31.port_b_first_address = 0;
defparam ram_block1a31.port_b_first_bit_number = 31;
defparam ram_block1a31.port_b_last_address = 31;
defparam ram_block1a31.port_b_logical_ram_depth = 32;
defparam ram_block1a31.port_b_logical_ram_width = 32;
defparam ram_block1a31.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a31.port_b_read_enable_clock = "clock0";
defparam ram_block1a31.ram_block_type = "auto";

cyclonev_ram_block ram_block1a21(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a21_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_register_bank_b_module:first_nios2_system_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_voi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a21.mixed_port_feed_through_mode = "old";
defparam ram_block1a21.operation_mode = "dual_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 5;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 31;
defparam ram_block1a21.port_a_logical_ram_depth = 32;
defparam ram_block1a21.port_a_logical_ram_width = 32;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a21.port_b_address_clear = "none";
defparam ram_block1a21.port_b_address_clock = "clock0";
defparam ram_block1a21.port_b_address_width = 5;
defparam ram_block1a21.port_b_data_out_clear = "none";
defparam ram_block1a21.port_b_data_out_clock = "none";
defparam ram_block1a21.port_b_data_width = 1;
defparam ram_block1a21.port_b_first_address = 0;
defparam ram_block1a21.port_b_first_bit_number = 21;
defparam ram_block1a21.port_b_last_address = 31;
defparam ram_block1a21.port_b_logical_ram_depth = 32;
defparam ram_block1a21.port_b_logical_ram_width = 32;
defparam ram_block1a21.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a21.port_b_read_enable_clock = "clock0";
defparam ram_block1a21.ram_block_type = "auto";

cyclonev_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_register_bank_b_module:first_nios2_system_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_voi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "old";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 5;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 31;
defparam ram_block1a11.port_a_logical_ram_depth = 32;
defparam ram_block1a11.port_a_logical_ram_width = 32;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock0";
defparam ram_block1a11.port_b_address_width = 5;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "none";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 31;
defparam ram_block1a11.port_b_logical_ram_depth = 32;
defparam ram_block1a11.port_b_logical_ram_width = 32;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock0";
defparam ram_block1a11.ram_block_type = "auto";

cyclonev_ram_block ram_block1a28(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[28]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a28_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a28.data_interleave_offset_in_bits = 1;
defparam ram_block1a28.data_interleave_width_in_bits = 1;
defparam ram_block1a28.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_register_bank_b_module:first_nios2_system_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_voi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a28.mixed_port_feed_through_mode = "old";
defparam ram_block1a28.operation_mode = "dual_port";
defparam ram_block1a28.port_a_address_clear = "none";
defparam ram_block1a28.port_a_address_width = 5;
defparam ram_block1a28.port_a_data_out_clear = "none";
defparam ram_block1a28.port_a_data_out_clock = "none";
defparam ram_block1a28.port_a_data_width = 1;
defparam ram_block1a28.port_a_first_address = 0;
defparam ram_block1a28.port_a_first_bit_number = 28;
defparam ram_block1a28.port_a_last_address = 31;
defparam ram_block1a28.port_a_logical_ram_depth = 32;
defparam ram_block1a28.port_a_logical_ram_width = 32;
defparam ram_block1a28.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a28.port_b_address_clear = "none";
defparam ram_block1a28.port_b_address_clock = "clock0";
defparam ram_block1a28.port_b_address_width = 5;
defparam ram_block1a28.port_b_data_out_clear = "none";
defparam ram_block1a28.port_b_data_out_clock = "none";
defparam ram_block1a28.port_b_data_width = 1;
defparam ram_block1a28.port_b_first_address = 0;
defparam ram_block1a28.port_b_first_bit_number = 28;
defparam ram_block1a28.port_b_last_address = 31;
defparam ram_block1a28.port_b_logical_ram_depth = 32;
defparam ram_block1a28.port_b_logical_ram_width = 32;
defparam ram_block1a28.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a28.port_b_read_enable_clock = "clock0";
defparam ram_block1a28.ram_block_type = "auto";

cyclonev_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_register_bank_b_module:first_nios2_system_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_voi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "old";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 5;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 31;
defparam ram_block1a10.port_a_logical_ram_depth = 32;
defparam ram_block1a10.port_a_logical_ram_width = 32;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock0";
defparam ram_block1a10.port_b_address_width = 5;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "none";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 31;
defparam ram_block1a10.port_b_logical_ram_depth = 32;
defparam ram_block1a10.port_b_logical_ram_width = 32;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock0";
defparam ram_block1a10.ram_block_type = "auto";

cyclonev_ram_block ram_block1a27(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[27]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a27_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a27.data_interleave_offset_in_bits = 1;
defparam ram_block1a27.data_interleave_width_in_bits = 1;
defparam ram_block1a27.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_register_bank_b_module:first_nios2_system_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_voi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a27.mixed_port_feed_through_mode = "old";
defparam ram_block1a27.operation_mode = "dual_port";
defparam ram_block1a27.port_a_address_clear = "none";
defparam ram_block1a27.port_a_address_width = 5;
defparam ram_block1a27.port_a_data_out_clear = "none";
defparam ram_block1a27.port_a_data_out_clock = "none";
defparam ram_block1a27.port_a_data_width = 1;
defparam ram_block1a27.port_a_first_address = 0;
defparam ram_block1a27.port_a_first_bit_number = 27;
defparam ram_block1a27.port_a_last_address = 31;
defparam ram_block1a27.port_a_logical_ram_depth = 32;
defparam ram_block1a27.port_a_logical_ram_width = 32;
defparam ram_block1a27.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a27.port_b_address_clear = "none";
defparam ram_block1a27.port_b_address_clock = "clock0";
defparam ram_block1a27.port_b_address_width = 5;
defparam ram_block1a27.port_b_data_out_clear = "none";
defparam ram_block1a27.port_b_data_out_clock = "none";
defparam ram_block1a27.port_b_data_width = 1;
defparam ram_block1a27.port_b_first_address = 0;
defparam ram_block1a27.port_b_first_bit_number = 27;
defparam ram_block1a27.port_b_last_address = 31;
defparam ram_block1a27.port_b_logical_ram_depth = 32;
defparam ram_block1a27.port_b_logical_ram_width = 32;
defparam ram_block1a27.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a27.port_b_read_enable_clock = "clock0";
defparam ram_block1a27.ram_block_type = "auto";

cyclonev_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_register_bank_b_module:first_nios2_system_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_voi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "old";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 5;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 31;
defparam ram_block1a8.port_a_logical_ram_depth = 32;
defparam ram_block1a8.port_a_logical_ram_width = 32;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock0";
defparam ram_block1a8.port_b_address_width = 5;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "none";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 31;
defparam ram_block1a8.port_b_logical_ram_depth = 32;
defparam ram_block1a8.port_b_logical_ram_width = 32;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock0";
defparam ram_block1a8.ram_block_type = "auto";

cyclonev_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_register_bank_b_module:first_nios2_system_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_voi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "old";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 5;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 31;
defparam ram_block1a9.port_a_logical_ram_depth = 32;
defparam ram_block1a9.port_a_logical_ram_width = 32;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock0";
defparam ram_block1a9.port_b_address_width = 5;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "none";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 31;
defparam ram_block1a9.port_b_logical_ram_depth = 32;
defparam ram_block1a9.port_b_logical_ram_width = 32;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock0";
defparam ram_block1a9.ram_block_type = "auto";

cyclonev_ram_block ram_block1a26(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[26]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a26_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a26.data_interleave_offset_in_bits = 1;
defparam ram_block1a26.data_interleave_width_in_bits = 1;
defparam ram_block1a26.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_register_bank_b_module:first_nios2_system_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_voi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a26.mixed_port_feed_through_mode = "old";
defparam ram_block1a26.operation_mode = "dual_port";
defparam ram_block1a26.port_a_address_clear = "none";
defparam ram_block1a26.port_a_address_width = 5;
defparam ram_block1a26.port_a_data_out_clear = "none";
defparam ram_block1a26.port_a_data_out_clock = "none";
defparam ram_block1a26.port_a_data_width = 1;
defparam ram_block1a26.port_a_first_address = 0;
defparam ram_block1a26.port_a_first_bit_number = 26;
defparam ram_block1a26.port_a_last_address = 31;
defparam ram_block1a26.port_a_logical_ram_depth = 32;
defparam ram_block1a26.port_a_logical_ram_width = 32;
defparam ram_block1a26.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a26.port_b_address_clear = "none";
defparam ram_block1a26.port_b_address_clock = "clock0";
defparam ram_block1a26.port_b_address_width = 5;
defparam ram_block1a26.port_b_data_out_clear = "none";
defparam ram_block1a26.port_b_data_out_clock = "none";
defparam ram_block1a26.port_b_data_width = 1;
defparam ram_block1a26.port_b_first_address = 0;
defparam ram_block1a26.port_b_first_bit_number = 26;
defparam ram_block1a26.port_b_last_address = 31;
defparam ram_block1a26.port_b_logical_ram_depth = 32;
defparam ram_block1a26.port_b_logical_ram_width = 32;
defparam ram_block1a26.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a26.port_b_read_enable_clock = "clock0";
defparam ram_block1a26.ram_block_type = "auto";

cyclonev_ram_block ram_block1a20(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a20_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_register_bank_b_module:first_nios2_system_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_voi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a20.mixed_port_feed_through_mode = "old";
defparam ram_block1a20.operation_mode = "dual_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 5;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 31;
defparam ram_block1a20.port_a_logical_ram_depth = 32;
defparam ram_block1a20.port_a_logical_ram_width = 32;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a20.port_b_address_clear = "none";
defparam ram_block1a20.port_b_address_clock = "clock0";
defparam ram_block1a20.port_b_address_width = 5;
defparam ram_block1a20.port_b_data_out_clear = "none";
defparam ram_block1a20.port_b_data_out_clock = "none";
defparam ram_block1a20.port_b_data_width = 1;
defparam ram_block1a20.port_b_first_address = 0;
defparam ram_block1a20.port_b_first_bit_number = 20;
defparam ram_block1a20.port_b_last_address = 31;
defparam ram_block1a20.port_b_logical_ram_depth = 32;
defparam ram_block1a20.port_b_logical_ram_width = 32;
defparam ram_block1a20.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a20.port_b_read_enable_clock = "clock0";
defparam ram_block1a20.ram_block_type = "auto";

cyclonev_ram_block ram_block1a19(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a19_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_register_bank_b_module:first_nios2_system_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_voi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a19.mixed_port_feed_through_mode = "old";
defparam ram_block1a19.operation_mode = "dual_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 5;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 31;
defparam ram_block1a19.port_a_logical_ram_depth = 32;
defparam ram_block1a19.port_a_logical_ram_width = 32;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a19.port_b_address_clear = "none";
defparam ram_block1a19.port_b_address_clock = "clock0";
defparam ram_block1a19.port_b_address_width = 5;
defparam ram_block1a19.port_b_data_out_clear = "none";
defparam ram_block1a19.port_b_data_out_clock = "none";
defparam ram_block1a19.port_b_data_width = 1;
defparam ram_block1a19.port_b_first_address = 0;
defparam ram_block1a19.port_b_first_bit_number = 19;
defparam ram_block1a19.port_b_last_address = 31;
defparam ram_block1a19.port_b_logical_ram_depth = 32;
defparam ram_block1a19.port_b_logical_ram_width = 32;
defparam ram_block1a19.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a19.port_b_read_enable_clock = "clock0";
defparam ram_block1a19.ram_block_type = "auto";

cyclonev_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_register_bank_b_module:first_nios2_system_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_voi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "old";
defparam ram_block1a17.operation_mode = "dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 5;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 31;
defparam ram_block1a17.port_a_logical_ram_depth = 32;
defparam ram_block1a17.port_a_logical_ram_width = 32;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a17.port_b_address_clear = "none";
defparam ram_block1a17.port_b_address_clock = "clock0";
defparam ram_block1a17.port_b_address_width = 5;
defparam ram_block1a17.port_b_data_out_clear = "none";
defparam ram_block1a17.port_b_data_out_clock = "none";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 31;
defparam ram_block1a17.port_b_logical_ram_depth = 32;
defparam ram_block1a17.port_b_logical_ram_width = 32;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock0";
defparam ram_block1a17.ram_block_type = "auto";

cyclonev_ram_block ram_block1a30(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[30]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a30_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a30.data_interleave_offset_in_bits = 1;
defparam ram_block1a30.data_interleave_width_in_bits = 1;
defparam ram_block1a30.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_register_bank_b_module:first_nios2_system_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_voi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a30.mixed_port_feed_through_mode = "old";
defparam ram_block1a30.operation_mode = "dual_port";
defparam ram_block1a30.port_a_address_clear = "none";
defparam ram_block1a30.port_a_address_width = 5;
defparam ram_block1a30.port_a_data_out_clear = "none";
defparam ram_block1a30.port_a_data_out_clock = "none";
defparam ram_block1a30.port_a_data_width = 1;
defparam ram_block1a30.port_a_first_address = 0;
defparam ram_block1a30.port_a_first_bit_number = 30;
defparam ram_block1a30.port_a_last_address = 31;
defparam ram_block1a30.port_a_logical_ram_depth = 32;
defparam ram_block1a30.port_a_logical_ram_width = 32;
defparam ram_block1a30.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a30.port_b_address_clear = "none";
defparam ram_block1a30.port_b_address_clock = "clock0";
defparam ram_block1a30.port_b_address_width = 5;
defparam ram_block1a30.port_b_data_out_clear = "none";
defparam ram_block1a30.port_b_data_out_clock = "none";
defparam ram_block1a30.port_b_data_width = 1;
defparam ram_block1a30.port_b_first_address = 0;
defparam ram_block1a30.port_b_first_bit_number = 30;
defparam ram_block1a30.port_b_last_address = 31;
defparam ram_block1a30.port_b_logical_ram_depth = 32;
defparam ram_block1a30.port_b_logical_ram_width = 32;
defparam ram_block1a30.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a30.port_b_read_enable_clock = "clock0";
defparam ram_block1a30.ram_block_type = "auto";

cyclonev_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_register_bank_b_module:first_nios2_system_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_voi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "old";
defparam ram_block1a18.operation_mode = "dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 5;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 31;
defparam ram_block1a18.port_a_logical_ram_depth = 32;
defparam ram_block1a18.port_a_logical_ram_width = 32;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a18.port_b_address_clear = "none";
defparam ram_block1a18.port_b_address_clock = "clock0";
defparam ram_block1a18.port_b_address_width = 5;
defparam ram_block1a18.port_b_data_out_clear = "none";
defparam ram_block1a18.port_b_data_out_clock = "none";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 31;
defparam ram_block1a18.port_b_logical_ram_depth = 32;
defparam ram_block1a18.port_b_logical_ram_width = 32;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock0";
defparam ram_block1a18.ram_block_type = "auto";

cyclonev_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_register_bank_b_module:first_nios2_system_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_voi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "old";
defparam ram_block1a16.operation_mode = "dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 5;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 31;
defparam ram_block1a16.port_a_logical_ram_depth = 32;
defparam ram_block1a16.port_a_logical_ram_width = 32;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a16.port_b_address_clear = "none";
defparam ram_block1a16.port_b_address_clock = "clock0";
defparam ram_block1a16.port_b_address_width = 5;
defparam ram_block1a16.port_b_data_out_clear = "none";
defparam ram_block1a16.port_b_data_out_clock = "none";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 31;
defparam ram_block1a16.port_b_logical_ram_depth = 32;
defparam ram_block1a16.port_b_logical_ram_width = 32;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock0";
defparam ram_block1a16.ram_block_type = "auto";

cyclonev_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_register_bank_b_module:first_nios2_system_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_voi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "old";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 5;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 31;
defparam ram_block1a15.port_a_logical_ram_depth = 32;
defparam ram_block1a15.port_a_logical_ram_width = 32;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock0";
defparam ram_block1a15.port_b_address_width = 5;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "none";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 31;
defparam ram_block1a15.port_b_logical_ram_depth = 32;
defparam ram_block1a15.port_b_logical_ram_width = 32;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock0";
defparam ram_block1a15.ram_block_type = "auto";

cyclonev_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_register_bank_b_module:first_nios2_system_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_voi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "old";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 5;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 31;
defparam ram_block1a12.port_a_logical_ram_depth = 32;
defparam ram_block1a12.port_a_logical_ram_width = 32;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock0";
defparam ram_block1a12.port_b_address_width = 5;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "none";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 31;
defparam ram_block1a12.port_b_logical_ram_depth = 32;
defparam ram_block1a12.port_b_logical_ram_width = 32;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock0";
defparam ram_block1a12.ram_block_type = "auto";

cyclonev_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_register_bank_b_module:first_nios2_system_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_voi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "old";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 5;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 31;
defparam ram_block1a13.port_a_logical_ram_depth = 32;
defparam ram_block1a13.port_a_logical_ram_width = 32;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock0";
defparam ram_block1a13.port_b_address_width = 5;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "none";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 31;
defparam ram_block1a13.port_b_logical_ram_depth = 32;
defparam ram_block1a13.port_b_logical_ram_width = 32;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock0";
defparam ram_block1a13.ram_block_type = "auto";

cyclonev_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_register_bank_b_module:first_nios2_system_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_voi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "old";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 5;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 31;
defparam ram_block1a14.port_a_logical_ram_depth = 32;
defparam ram_block1a14.port_a_logical_ram_width = 32;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock0";
defparam ram_block1a14.port_b_address_width = 5;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "none";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 31;
defparam ram_block1a14.port_b_logical_ram_depth = 32;
defparam ram_block1a14.port_b_logical_ram_width = 32;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock0";
defparam ram_block1a14.ram_block_type = "auto";

cyclonev_ram_block ram_block1a29(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[29]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a29_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a29.data_interleave_offset_in_bits = 1;
defparam ram_block1a29.data_interleave_width_in_bits = 1;
defparam ram_block1a29.logical_ram_name = "first_nios2_system_cpu:cpu|first_nios2_system_cpu_cpu:cpu|first_nios2_system_cpu_cpu_register_bank_b_module:first_nios2_system_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_voi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a29.mixed_port_feed_through_mode = "old";
defparam ram_block1a29.operation_mode = "dual_port";
defparam ram_block1a29.port_a_address_clear = "none";
defparam ram_block1a29.port_a_address_width = 5;
defparam ram_block1a29.port_a_data_out_clear = "none";
defparam ram_block1a29.port_a_data_out_clock = "none";
defparam ram_block1a29.port_a_data_width = 1;
defparam ram_block1a29.port_a_first_address = 0;
defparam ram_block1a29.port_a_first_bit_number = 29;
defparam ram_block1a29.port_a_last_address = 31;
defparam ram_block1a29.port_a_logical_ram_depth = 32;
defparam ram_block1a29.port_a_logical_ram_width = 32;
defparam ram_block1a29.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a29.port_b_address_clear = "none";
defparam ram_block1a29.port_b_address_clock = "clock0";
defparam ram_block1a29.port_b_address_width = 5;
defparam ram_block1a29.port_b_data_out_clear = "none";
defparam ram_block1a29.port_b_data_out_clock = "none";
defparam ram_block1a29.port_b_data_width = 1;
defparam ram_block1a29.port_b_first_address = 0;
defparam ram_block1a29.port_b_first_bit_number = 29;
defparam ram_block1a29.port_b_last_address = 31;
defparam ram_block1a29.port_b_logical_ram_depth = 32;
defparam ram_block1a29.port_b_logical_ram_width = 32;
defparam ram_block1a29.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a29.port_b_read_enable_clock = "clock0";
defparam ram_block1a29.ram_block_type = "auto";

endmodule

module first_nios2_system_first_nios2_system_download1 (
	data_out1,
	A_st_data_0,
	mem_used_1,
	Equal15,
	always0,
	clr_break_line,
	wait_latency_counter_1,
	wait_latency_counter_0,
	d_write,
	Equal0,
	reset_n,
	clk)/* synthesis synthesis_greybox=1 */;
output 	data_out1;
input 	A_st_data_0;
input 	mem_used_1;
input 	Equal15;
output 	always0;
input 	clr_break_line;
input 	wait_latency_counter_1;
input 	wait_latency_counter_0;
input 	d_write;
input 	Equal0;
input 	reset_n;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \always0~1_combout ;
wire \data_out~0_combout ;


dffeas data_out(
	.clk(clk),
	.d(\data_out~0_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out1),
	.prn(vcc));
defparam data_out.is_wysiwyg = "true";
defparam data_out.power_up = "low";

cyclonev_lcell_comb \always0~0 (
	.dataa(!mem_used_1),
	.datab(!Equal15),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(always0),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \always0~0 .shared_arith = "off";

cyclonev_lcell_comb \always0~1 (
	.dataa(!clr_break_line),
	.datab(!wait_latency_counter_1),
	.datac(!wait_latency_counter_0),
	.datad(!d_write),
	.datae(!Equal0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~1 .extended_lut = "off";
defparam \always0~1 .lut_mask = 64'hFFFFFDFFFFFFFDFF;
defparam \always0~1 .shared_arith = "off";

cyclonev_lcell_comb \data_out~0 (
	.dataa(!data_out1),
	.datab(!A_st_data_0),
	.datac(!always0),
	.datad(!\always0~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~0 .extended_lut = "off";
defparam \data_out~0 .lut_mask = 64'h7FF77FF77FF77FF7;
defparam \data_out~0 .shared_arith = "off";

endmodule

module first_nios2_system_first_nios2_system_download1_1 (
	data_out1,
	A_st_data_0,
	clr_break_line,
	d_write,
	Equal0,
	reset_n,
	write,
	wait_latency_counter_0,
	clk)/* synthesis synthesis_greybox=1 */;
output 	data_out1;
input 	A_st_data_0;
input 	clr_break_line;
input 	d_write;
input 	Equal0;
input 	reset_n;
input 	write;
input 	wait_latency_counter_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \always0~0_combout ;
wire \data_out~0_combout ;


dffeas data_out(
	.clk(clk),
	.d(\data_out~0_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out1),
	.prn(vcc));
defparam data_out.is_wysiwyg = "true";
defparam data_out.power_up = "low";

cyclonev_lcell_comb \always0~0 (
	.dataa(!d_write),
	.datab(!Equal0),
	.datac(!wait_latency_counter_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'hFDFDFDFDFDFDFDFD;
defparam \always0~0 .shared_arith = "off";

cyclonev_lcell_comb \data_out~0 (
	.dataa(!data_out1),
	.datab(!A_st_data_0),
	.datac(!clr_break_line),
	.datad(!write),
	.datae(!\always0~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~0 .extended_lut = "off";
defparam \data_out~0 .lut_mask = 64'hF77F7FF7F77F7FF7;
defparam \data_out~0 .shared_arith = "off";

endmodule

module first_nios2_system_first_nios2_system_download1_2 (
	data_out1,
	A_st_data_0,
	clr_break_line,
	d_write,
	Equal0,
	reset_n,
	wait_latency_counter_1,
	m0_write,
	wait_latency_counter_0,
	clk)/* synthesis synthesis_greybox=1 */;
output 	data_out1;
input 	A_st_data_0;
input 	clr_break_line;
input 	d_write;
input 	Equal0;
input 	reset_n;
input 	wait_latency_counter_1;
input 	m0_write;
input 	wait_latency_counter_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \always0~0_combout ;
wire \data_out~0_combout ;


dffeas data_out(
	.clk(clk),
	.d(\data_out~0_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out1),
	.prn(vcc));
defparam data_out.is_wysiwyg = "true";
defparam data_out.power_up = "low";

cyclonev_lcell_comb \always0~0 (
	.dataa(!d_write),
	.datab(!Equal0),
	.datac(!wait_latency_counter_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'hFDFDFDFDFDFDFDFD;
defparam \always0~0 .shared_arith = "off";

cyclonev_lcell_comb \data_out~0 (
	.dataa(!data_out1),
	.datab(!A_st_data_0),
	.datac(!clr_break_line),
	.datad(!wait_latency_counter_1),
	.datae(!m0_write),
	.dataf(!\always0~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~0 .extended_lut = "off";
defparam \data_out~0 .lut_mask = 64'h7FF7F77FF77F7FF7;
defparam \data_out~0 .shared_arith = "off";

endmodule

module first_nios2_system_first_nios2_system_hex1 (
	data_out_0,
	data_out_1,
	data_out_2,
	data_out_3,
	data_out_4,
	data_out_5,
	data_out_6,
	writedata,
	clr_break_line,
	d_write,
	Equal0,
	reset_n,
	wait_latency_counter_1,
	mem_used_1,
	Equal6,
	wait_latency_counter_0,
	clk)/* synthesis synthesis_greybox=1 */;
output 	data_out_0;
output 	data_out_1;
output 	data_out_2;
output 	data_out_3;
output 	data_out_4;
output 	data_out_5;
output 	data_out_6;
input 	[31:0] writedata;
input 	clr_break_line;
input 	d_write;
input 	Equal0;
input 	reset_n;
input 	wait_latency_counter_1;
input 	mem_used_1;
input 	Equal6;
input 	wait_latency_counter_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \always0~0_combout ;
wire \always0~1_combout ;


dffeas \data_out[0] (
	.clk(clk),
	.d(writedata[0]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_0),
	.prn(vcc));
defparam \data_out[0] .is_wysiwyg = "true";
defparam \data_out[0] .power_up = "low";

dffeas \data_out[1] (
	.clk(clk),
	.d(writedata[1]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_1),
	.prn(vcc));
defparam \data_out[1] .is_wysiwyg = "true";
defparam \data_out[1] .power_up = "low";

dffeas \data_out[2] (
	.clk(clk),
	.d(writedata[2]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_2),
	.prn(vcc));
defparam \data_out[2] .is_wysiwyg = "true";
defparam \data_out[2] .power_up = "low";

dffeas \data_out[3] (
	.clk(clk),
	.d(writedata[3]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_3),
	.prn(vcc));
defparam \data_out[3] .is_wysiwyg = "true";
defparam \data_out[3] .power_up = "low";

dffeas \data_out[4] (
	.clk(clk),
	.d(writedata[4]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_4),
	.prn(vcc));
defparam \data_out[4] .is_wysiwyg = "true";
defparam \data_out[4] .power_up = "low";

dffeas \data_out[5] (
	.clk(clk),
	.d(writedata[5]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_5),
	.prn(vcc));
defparam \data_out[5] .is_wysiwyg = "true";
defparam \data_out[5] .power_up = "low";

dffeas \data_out[6] (
	.clk(clk),
	.d(writedata[6]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_6),
	.prn(vcc));
defparam \data_out[6] .is_wysiwyg = "true";
defparam \data_out[6] .power_up = "low";

cyclonev_lcell_comb \always0~0 (
	.dataa(!d_write),
	.datab(!Equal0),
	.datac(!wait_latency_counter_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'hFDFDFDFDFDFDFDFD;
defparam \always0~0 .shared_arith = "off";

cyclonev_lcell_comb \always0~1 (
	.dataa(!clr_break_line),
	.datab(!wait_latency_counter_1),
	.datac(!mem_used_1),
	.datad(!Equal6),
	.datae(!\always0~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~1 .extended_lut = "off";
defparam \always0~1 .lut_mask = 64'hFDFFFFFFFDFFFFFF;
defparam \always0~1 .shared_arith = "off";

endmodule

module first_nios2_system_first_nios2_system_hex1_1 (
	data_out_0,
	data_out_1,
	data_out_2,
	data_out_3,
	data_out_4,
	data_out_5,
	data_out_6,
	writedata,
	A_mem_baddr_7,
	clr_break_line,
	d_write,
	Equal0,
	reset_n,
	wait_latency_counter_1,
	mem_used_1,
	always1,
	wait_latency_counter_0,
	clk)/* synthesis synthesis_greybox=1 */;
output 	data_out_0;
output 	data_out_1;
output 	data_out_2;
output 	data_out_3;
output 	data_out_4;
output 	data_out_5;
output 	data_out_6;
input 	[31:0] writedata;
input 	A_mem_baddr_7;
input 	clr_break_line;
input 	d_write;
input 	Equal0;
input 	reset_n;
input 	wait_latency_counter_1;
input 	mem_used_1;
input 	always1;
input 	wait_latency_counter_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \always0~0_combout ;
wire \always0~1_combout ;


dffeas \data_out[0] (
	.clk(clk),
	.d(writedata[0]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_0),
	.prn(vcc));
defparam \data_out[0] .is_wysiwyg = "true";
defparam \data_out[0] .power_up = "low";

dffeas \data_out[1] (
	.clk(clk),
	.d(writedata[1]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_1),
	.prn(vcc));
defparam \data_out[1] .is_wysiwyg = "true";
defparam \data_out[1] .power_up = "low";

dffeas \data_out[2] (
	.clk(clk),
	.d(writedata[2]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_2),
	.prn(vcc));
defparam \data_out[2] .is_wysiwyg = "true";
defparam \data_out[2] .power_up = "low";

dffeas \data_out[3] (
	.clk(clk),
	.d(writedata[3]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_3),
	.prn(vcc));
defparam \data_out[3] .is_wysiwyg = "true";
defparam \data_out[3] .power_up = "low";

dffeas \data_out[4] (
	.clk(clk),
	.d(writedata[4]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_4),
	.prn(vcc));
defparam \data_out[4] .is_wysiwyg = "true";
defparam \data_out[4] .power_up = "low";

dffeas \data_out[5] (
	.clk(clk),
	.d(writedata[5]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_5),
	.prn(vcc));
defparam \data_out[5] .is_wysiwyg = "true";
defparam \data_out[5] .power_up = "low";

dffeas \data_out[6] (
	.clk(clk),
	.d(writedata[6]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_6),
	.prn(vcc));
defparam \data_out[6] .is_wysiwyg = "true";
defparam \data_out[6] .power_up = "low";

cyclonev_lcell_comb \always0~0 (
	.dataa(!d_write),
	.datab(!Equal0),
	.datac(!wait_latency_counter_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'hFDFDFDFDFDFDFDFD;
defparam \always0~0 .shared_arith = "off";

cyclonev_lcell_comb \always0~1 (
	.dataa(!clr_break_line),
	.datab(!A_mem_baddr_7),
	.datac(!wait_latency_counter_1),
	.datad(!mem_used_1),
	.datae(!always1),
	.dataf(!\always0~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~1 .extended_lut = "off";
defparam \always0~1 .lut_mask = 64'hFFFDFFFFFFFFFFFF;
defparam \always0~1 .shared_arith = "off";

endmodule

module first_nios2_system_first_nios2_system_jtag_uart (
	q_b_0,
	q_b_1,
	q_b_2,
	q_b_3,
	q_b_4,
	q_b_5,
	q_b_6,
	q_b_7,
	Add1,
	Add11,
	Add12,
	Add13,
	Add14,
	Add15,
	Add16,
	tdo,
	A_st_data_0,
	A_mem_baddr_4,
	Equal1,
	Equal2,
	clr_break_line,
	d_write,
	A_mem_baddr_3,
	A_mem_baddr_2,
	r_sync_rst,
	A_st_data_1,
	A_st_data_2,
	A_st_data_3,
	A_st_data_4,
	A_st_data_5,
	A_st_data_6,
	A_st_data_7,
	read_latency_shift_reg,
	cp_valid,
	always1,
	av_waitrequest1,
	mem_used_1,
	av_waitrequest2,
	ien_AE1,
	av_readdata_9,
	ien_AF1,
	av_readdata_8,
	b_full,
	b_full1,
	b_non_empty,
	read_01,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_5,
	A_st_data_10,
	ac1,
	rvalid1,
	woverflow1,
	altera_internal_jtag,
	altera_internal_jtag1,
	state_4,
	splitter_nodes_receive_0_3,
	virtual_ir_scan_reg,
	clr_reg,
	state_3,
	state_8,
	irf_reg_0_1,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_0;
output 	q_b_1;
output 	q_b_2;
output 	q_b_3;
output 	q_b_4;
output 	q_b_5;
output 	q_b_6;
output 	q_b_7;
output 	Add1;
output 	Add11;
output 	Add12;
output 	Add13;
output 	Add14;
output 	Add15;
output 	Add16;
output 	tdo;
input 	A_st_data_0;
input 	A_mem_baddr_4;
input 	Equal1;
input 	Equal2;
input 	clr_break_line;
input 	d_write;
input 	A_mem_baddr_3;
input 	A_mem_baddr_2;
input 	r_sync_rst;
input 	A_st_data_1;
input 	A_st_data_2;
input 	A_st_data_3;
input 	A_st_data_4;
input 	A_st_data_5;
input 	A_st_data_6;
input 	A_st_data_7;
input 	read_latency_shift_reg;
input 	cp_valid;
input 	always1;
output 	av_waitrequest1;
input 	mem_used_1;
output 	av_waitrequest2;
output 	ien_AE1;
output 	av_readdata_9;
output 	ien_AF1;
output 	av_readdata_8;
output 	b_full;
output 	b_full1;
output 	b_non_empty;
output 	read_01;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_5;
input 	A_st_data_10;
output 	ac1;
output 	rvalid1;
output 	woverflow1;
input 	altera_internal_jtag;
input 	altera_internal_jtag1;
input 	state_4;
input 	splitter_nodes_receive_0_3;
input 	virtual_ir_scan_reg;
input 	clr_reg;
input 	state_3;
input 	state_8;
input 	irf_reg_0_1;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \the_first_nios2_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[7] ;
wire \the_first_nios2_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[0] ;
wire \the_first_nios2_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[1] ;
wire \the_first_nios2_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[2] ;
wire \the_first_nios2_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[3] ;
wire \the_first_nios2_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[4] ;
wire \the_first_nios2_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[5] ;
wire \the_first_nios2_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[6] ;
wire \t_dav~q ;
wire \r_val~q ;
wire \the_first_nios2_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[3]~q ;
wire \the_first_nios2_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[0]~q ;
wire \the_first_nios2_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[2]~q ;
wire \the_first_nios2_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[1]~q ;
wire \the_first_nios2_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[5]~q ;
wire \the_first_nios2_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[4]~q ;
wire \first_nios2_system_jtag_uart_alt_jtag_atlantic|t_pause~q ;
wire \fifo_wr~q ;
wire \first_nios2_system_jtag_uart_alt_jtag_atlantic|rvalid0~1_combout ;
wire \the_first_nios2_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|b_non_empty~q ;
wire \r_val~0_combout ;
wire \fifo_rd~0_combout ;
wire \first_nios2_system_jtag_uart_alt_jtag_atlantic|t_ena~q ;
wire \wr_rfifo~combout ;
wire \fifo_wr~0_combout ;
wire \first_nios2_system_jtag_uart_alt_jtag_atlantic|wdata[0]~q ;
wire \first_nios2_system_jtag_uart_alt_jtag_atlantic|wdata[1]~q ;
wire \first_nios2_system_jtag_uart_alt_jtag_atlantic|wdata[2]~q ;
wire \first_nios2_system_jtag_uart_alt_jtag_atlantic|wdata[3]~q ;
wire \first_nios2_system_jtag_uart_alt_jtag_atlantic|wdata[4]~q ;
wire \first_nios2_system_jtag_uart_alt_jtag_atlantic|wdata[5]~q ;
wire \first_nios2_system_jtag_uart_alt_jtag_atlantic|wdata[6]~q ;
wire \first_nios2_system_jtag_uart_alt_jtag_atlantic|wdata[7]~q ;
wire \Add1~6 ;
wire \Add1~10 ;
wire \Add1~14 ;
wire \Add1~18 ;
wire \Add1~22 ;
wire \Add1~26 ;
wire \av_waitrequest~1_combout ;
wire \ien_AE~0_combout ;
wire \LessThan0~0_combout ;
wire \LessThan0~1_combout ;
wire \fifo_AE~q ;
wire \pause_irq~0_combout ;
wire \pause_irq~q ;
wire \Add0~22 ;
wire \Add0~26 ;
wire \Add0~18 ;
wire \Add0~1_sumout ;
wire \Add0~2 ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \Add0~13_sumout ;
wire \Add0~17_sumout ;
wire \Add0~21_sumout ;
wire \Add0~25_sumout ;
wire \LessThan1~0_combout ;
wire \LessThan1~1_combout ;
wire \fifo_AF~q ;
wire \fifo_rd~1_combout ;
wire \ac~0_combout ;
wire \rvalid~0_combout ;
wire \woverflow~0_combout ;
wire \woverflow~1_combout ;


first_nios2_system_alt_jtag_atlantic first_nios2_system_jtag_uart_alt_jtag_atlantic(
	.r_dat({\the_first_nios2_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[7] ,\the_first_nios2_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[6] ,
\the_first_nios2_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[5] ,\the_first_nios2_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[4] ,
\the_first_nios2_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[3] ,\the_first_nios2_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[2] ,
\the_first_nios2_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[1] ,\the_first_nios2_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[0] }),
	.tdo1(tdo),
	.clr_break_line(clr_break_line),
	.rst_n(r_sync_rst),
	.t_dav(\t_dav~q ),
	.r_val(\r_val~q ),
	.t_pause1(\first_nios2_system_jtag_uart_alt_jtag_atlantic|t_pause~q ),
	.rvalid01(\first_nios2_system_jtag_uart_alt_jtag_atlantic|rvalid0~1_combout ),
	.t_ena1(\first_nios2_system_jtag_uart_alt_jtag_atlantic|t_ena~q ),
	.wdata_0(\first_nios2_system_jtag_uart_alt_jtag_atlantic|wdata[0]~q ),
	.wdata_1(\first_nios2_system_jtag_uart_alt_jtag_atlantic|wdata[1]~q ),
	.wdata_2(\first_nios2_system_jtag_uart_alt_jtag_atlantic|wdata[2]~q ),
	.wdata_3(\first_nios2_system_jtag_uart_alt_jtag_atlantic|wdata[3]~q ),
	.wdata_4(\first_nios2_system_jtag_uart_alt_jtag_atlantic|wdata[4]~q ),
	.wdata_5(\first_nios2_system_jtag_uart_alt_jtag_atlantic|wdata[5]~q ),
	.wdata_6(\first_nios2_system_jtag_uart_alt_jtag_atlantic|wdata[6]~q ),
	.wdata_7(\first_nios2_system_jtag_uart_alt_jtag_atlantic|wdata[7]~q ),
	.altera_internal_jtag(altera_internal_jtag),
	.altera_internal_jtag1(altera_internal_jtag1),
	.state_4(state_4),
	.splitter_nodes_receive_0_3(splitter_nodes_receive_0_3),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.clr_reg(clr_reg),
	.state_3(state_3),
	.state_8(state_8),
	.irf_reg_0_1(irf_reg_0_1),
	.clk(clk_clk));

first_nios2_system_first_nios2_system_jtag_uart_scfifo_r the_first_nios2_system_jtag_uart_scfifo_r(
	.q_b_0(q_b_0),
	.q_b_1(q_b_1),
	.q_b_2(q_b_2),
	.q_b_3(q_b_3),
	.q_b_4(q_b_4),
	.q_b_5(q_b_5),
	.q_b_6(q_b_6),
	.q_b_7(q_b_7),
	.A_mem_baddr_2(A_mem_baddr_2),
	.r_sync_rst(r_sync_rst),
	.read_latency_shift_reg(read_latency_shift_reg),
	.av_waitrequest(av_waitrequest1),
	.av_waitrequest1(av_waitrequest2),
	.b_full(b_full),
	.b_non_empty(b_non_empty),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_1(counter_reg_bit_1),
	.fifo_rd(\fifo_rd~0_combout ),
	.t_ena(\first_nios2_system_jtag_uart_alt_jtag_atlantic|t_ena~q ),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_5(counter_reg_bit_5),
	.wr_rfifo(\wr_rfifo~combout ),
	.wdata_0(\first_nios2_system_jtag_uart_alt_jtag_atlantic|wdata[0]~q ),
	.wdata_1(\first_nios2_system_jtag_uart_alt_jtag_atlantic|wdata[1]~q ),
	.wdata_2(\first_nios2_system_jtag_uart_alt_jtag_atlantic|wdata[2]~q ),
	.wdata_3(\first_nios2_system_jtag_uart_alt_jtag_atlantic|wdata[3]~q ),
	.wdata_4(\first_nios2_system_jtag_uart_alt_jtag_atlantic|wdata[4]~q ),
	.wdata_5(\first_nios2_system_jtag_uart_alt_jtag_atlantic|wdata[5]~q ),
	.wdata_6(\first_nios2_system_jtag_uart_alt_jtag_atlantic|wdata[6]~q ),
	.wdata_7(\first_nios2_system_jtag_uart_alt_jtag_atlantic|wdata[7]~q ),
	.clk_clk(clk_clk));

first_nios2_system_first_nios2_system_jtag_uart_scfifo_w the_first_nios2_system_jtag_uart_scfifo_w(
	.q_b_7(\the_first_nios2_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.q_b_0(\the_first_nios2_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[0] ),
	.q_b_1(\the_first_nios2_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[1] ),
	.q_b_2(\the_first_nios2_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[2] ),
	.q_b_3(\the_first_nios2_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[3] ),
	.q_b_4(\the_first_nios2_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[4] ),
	.q_b_5(\the_first_nios2_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.q_b_6(\the_first_nios2_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.A_st_data_0(A_st_data_0),
	.r_sync_rst(r_sync_rst),
	.A_st_data_1(A_st_data_1),
	.A_st_data_2(A_st_data_2),
	.A_st_data_3(A_st_data_3),
	.A_st_data_4(A_st_data_4),
	.A_st_data_5(A_st_data_5),
	.A_st_data_6(A_st_data_6),
	.A_st_data_7(A_st_data_7),
	.b_full(b_full1),
	.counter_reg_bit_3(\the_first_nios2_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[3]~q ),
	.counter_reg_bit_0(\the_first_nios2_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[0]~q ),
	.counter_reg_bit_2(\the_first_nios2_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[2]~q ),
	.counter_reg_bit_1(\the_first_nios2_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[1]~q ),
	.counter_reg_bit_5(\the_first_nios2_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[5]~q ),
	.counter_reg_bit_4(\the_first_nios2_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[4]~q ),
	.fifo_wr(\fifo_wr~q ),
	.rvalid0(\first_nios2_system_jtag_uart_alt_jtag_atlantic|rvalid0~1_combout ),
	.b_non_empty(\the_first_nios2_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|b_non_empty~q ),
	.r_val(\r_val~0_combout ),
	.clk_clk(clk_clk));

dffeas t_dav(
	.clk(clk_clk),
	.d(b_full),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\t_dav~q ),
	.prn(vcc));
defparam t_dav.is_wysiwyg = "true";
defparam t_dav.power_up = "low";

dffeas r_val(
	.clk(clk_clk),
	.d(\r_val~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\r_val~q ),
	.prn(vcc));
defparam r_val.is_wysiwyg = "true";
defparam r_val.power_up = "low";

dffeas fifo_wr(
	.clk(clk_clk),
	.d(\fifo_wr~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\fifo_wr~q ),
	.prn(vcc));
defparam fifo_wr.is_wysiwyg = "true";
defparam fifo_wr.power_up = "low";

cyclonev_lcell_comb \r_val~0 (
	.dataa(!\first_nios2_system_jtag_uart_alt_jtag_atlantic|rvalid0~1_combout ),
	.datab(!\the_first_nios2_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|b_non_empty~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\r_val~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \r_val~0 .extended_lut = "off";
defparam \r_val~0 .lut_mask = 64'h7777777777777777;
defparam \r_val~0 .shared_arith = "off";

cyclonev_lcell_comb \fifo_rd~0 (
	.dataa(!A_mem_baddr_2),
	.datab(!av_waitrequest1),
	.datac(!av_waitrequest2),
	.datad(!read_latency_shift_reg),
	.datae(!b_non_empty),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fifo_rd~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_rd~0 .extended_lut = "off";
defparam \fifo_rd~0 .lut_mask = 64'hEFFFFFFFEFFFFFFF;
defparam \fifo_rd~0 .shared_arith = "off";

cyclonev_lcell_comb wr_rfifo(
	.dataa(!b_full),
	.datab(!\first_nios2_system_jtag_uart_alt_jtag_atlantic|t_ena~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wr_rfifo~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam wr_rfifo.extended_lut = "off";
defparam wr_rfifo.lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam wr_rfifo.shared_arith = "off";

cyclonev_lcell_comb \fifo_wr~0 (
	.dataa(!b_full1),
	.datab(!\woverflow~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fifo_wr~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_wr~0 .extended_lut = "off";
defparam \fifo_wr~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \fifo_wr~0 .shared_arith = "off";

cyclonev_lcell_comb \Add1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!b_full1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add1),
	.cout(),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h000000000000FF00;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \Add1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\the_first_nios2_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add11),
	.cout(\Add1~6 ),
	.shareout());
defparam \Add1~5 .extended_lut = "off";
defparam \Add1~5 .lut_mask = 64'h000000000000FF00;
defparam \Add1~5 .shared_arith = "off";

cyclonev_lcell_comb \Add1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\the_first_nios2_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add12),
	.cout(\Add1~10 ),
	.shareout());
defparam \Add1~9 .extended_lut = "off";
defparam \Add1~9 .lut_mask = 64'h000000000000FF00;
defparam \Add1~9 .shared_arith = "off";

cyclonev_lcell_comb \Add1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\the_first_nios2_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add13),
	.cout(\Add1~14 ),
	.shareout());
defparam \Add1~13 .extended_lut = "off";
defparam \Add1~13 .lut_mask = 64'h000000000000FF00;
defparam \Add1~13 .shared_arith = "off";

cyclonev_lcell_comb \Add1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\the_first_nios2_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add14),
	.cout(\Add1~18 ),
	.shareout());
defparam \Add1~17 .extended_lut = "off";
defparam \Add1~17 .lut_mask = 64'h000000000000FF00;
defparam \Add1~17 .shared_arith = "off";

cyclonev_lcell_comb \Add1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\the_first_nios2_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add15),
	.cout(\Add1~22 ),
	.shareout());
defparam \Add1~21 .extended_lut = "off";
defparam \Add1~21 .lut_mask = 64'h000000000000FF00;
defparam \Add1~21 .shared_arith = "off";

cyclonev_lcell_comb \Add1~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\the_first_nios2_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Add16),
	.cout(\Add1~26 ),
	.shareout());
defparam \Add1~25 .extended_lut = "off";
defparam \Add1~25 .lut_mask = 64'h000000000000FF00;
defparam \Add1~25 .shared_arith = "off";

dffeas av_waitrequest(
	.clk(clk_clk),
	.d(\av_waitrequest~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_waitrequest1),
	.prn(vcc));
defparam av_waitrequest.is_wysiwyg = "true";
defparam av_waitrequest.power_up = "low";

cyclonev_lcell_comb \av_waitrequest~0 (
	.dataa(!A_mem_baddr_3),
	.datab(!A_mem_baddr_4),
	.datac(!Equal1),
	.datad(!Equal2),
	.datae(!mem_used_1),
	.dataf(!always1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(av_waitrequest2),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_waitrequest~0 .extended_lut = "off";
defparam \av_waitrequest~0 .lut_mask = 64'hFFFFDFFFFFFFFFFF;
defparam \av_waitrequest~0 .shared_arith = "off";

dffeas ien_AE(
	.clk(clk_clk),
	.d(A_st_data_1),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ien_AE~0_combout ),
	.q(ien_AE1),
	.prn(vcc));
defparam ien_AE.is_wysiwyg = "true";
defparam ien_AE.power_up = "low";

cyclonev_lcell_comb \av_readdata[9] (
	.dataa(!\fifo_AE~q ),
	.datab(!ien_AE1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(av_readdata_9),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_readdata[9] .extended_lut = "off";
defparam \av_readdata[9] .lut_mask = 64'h7777777777777777;
defparam \av_readdata[9] .shared_arith = "off";

dffeas ien_AF(
	.clk(clk_clk),
	.d(A_st_data_0),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ien_AE~0_combout ),
	.q(ien_AF1),
	.prn(vcc));
defparam ien_AF.is_wysiwyg = "true";
defparam ien_AF.power_up = "low";

cyclonev_lcell_comb \av_readdata[8]~0 (
	.dataa(!ien_AF1),
	.datab(!\pause_irq~q ),
	.datac(!\fifo_AF~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(av_readdata_8),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_readdata[8]~0 .extended_lut = "off";
defparam \av_readdata[8]~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \av_readdata[8]~0 .shared_arith = "off";

dffeas read_0(
	.clk(clk_clk),
	.d(\fifo_rd~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_01),
	.prn(vcc));
defparam read_0.is_wysiwyg = "true";
defparam read_0.power_up = "low";

dffeas ac(
	.clk(clk_clk),
	.d(\ac~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ac1),
	.prn(vcc));
defparam ac.is_wysiwyg = "true";
defparam ac.power_up = "low";

dffeas rvalid(
	.clk(clk_clk),
	.d(\rvalid~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(rvalid1),
	.prn(vcc));
defparam rvalid.is_wysiwyg = "true";
defparam rvalid.power_up = "low";

dffeas woverflow(
	.clk(clk_clk),
	.d(\woverflow~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(woverflow1),
	.prn(vcc));
defparam woverflow.is_wysiwyg = "true";
defparam woverflow.power_up = "low";

cyclonev_lcell_comb \av_waitrequest~1 (
	.dataa(!cp_valid),
	.datab(!av_waitrequest1),
	.datac(!av_waitrequest2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_waitrequest~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_waitrequest~1 .extended_lut = "off";
defparam \av_waitrequest~1 .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \av_waitrequest~1 .shared_arith = "off";

cyclonev_lcell_comb \ien_AE~0 (
	.dataa(!clr_break_line),
	.datab(!d_write),
	.datac(!A_mem_baddr_2),
	.datad(!av_waitrequest1),
	.datae(!av_waitrequest2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ien_AE~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ien_AE~0 .extended_lut = "off";
defparam \ien_AE~0 .lut_mask = 64'hFF7FFFFFFF7FFFFF;
defparam \ien_AE~0 .shared_arith = "off";

cyclonev_lcell_comb \LessThan0~0 (
	.dataa(!\the_first_nios2_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[3]~q ),
	.datab(!\the_first_nios2_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[0]~q ),
	.datac(!\the_first_nios2_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[2]~q ),
	.datad(!\the_first_nios2_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~0 .extended_lut = "off";
defparam \LessThan0~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \LessThan0~0 .shared_arith = "off";

cyclonev_lcell_comb \LessThan0~1 (
	.dataa(!b_full1),
	.datab(!\LessThan0~0_combout ),
	.datac(!\the_first_nios2_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[5]~q ),
	.datad(!\the_first_nios2_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~1 .extended_lut = "off";
defparam \LessThan0~1 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \LessThan0~1 .shared_arith = "off";

dffeas fifo_AE(
	.clk(clk_clk),
	.d(\LessThan0~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\fifo_AE~q ),
	.prn(vcc));
defparam fifo_AE.is_wysiwyg = "true";
defparam fifo_AE.power_up = "low";

cyclonev_lcell_comb \pause_irq~0 (
	.dataa(!\pause_irq~q ),
	.datab(!b_non_empty),
	.datac(!\first_nios2_system_jtag_uart_alt_jtag_atlantic|t_pause~q ),
	.datad(!read_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pause_irq~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pause_irq~0 .extended_lut = "off";
defparam \pause_irq~0 .lut_mask = 64'hFF7FFF7FFF7FFF7F;
defparam \pause_irq~0 .shared_arith = "off";

dffeas pause_irq(
	.clk(clk_clk),
	.d(\pause_irq~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\pause_irq~q ),
	.prn(vcc));
defparam pause_irq.is_wysiwyg = "true";
defparam pause_irq.power_up = "low";

cyclonev_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_0),
	.datae(gnd),
	.dataf(!counter_reg_bit_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~21 .shared_arith = "off";

cyclonev_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h000000000000FF00;
defparam \Add0~25 .shared_arith = "off";

cyclonev_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h000000000000FF00;
defparam \Add0~17 .shared_arith = "off";

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(\Add0~2 ),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h000000000000FF00;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h000000000000FF00;
defparam \Add0~5 .shared_arith = "off";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!b_full),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h000000000000FF00;
defparam \Add0~9 .shared_arith = "off";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000000000000000;
defparam \Add0~13 .shared_arith = "off";

cyclonev_lcell_comb \LessThan1~0 (
	.dataa(!counter_reg_bit_0),
	.datab(!\Add0~17_sumout ),
	.datac(!\Add0~21_sumout ),
	.datad(!\Add0~25_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan1~0 .extended_lut = "off";
defparam \LessThan1~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \LessThan1~0 .shared_arith = "off";

cyclonev_lcell_comb \LessThan1~1 (
	.dataa(!\Add0~1_sumout ),
	.datab(!\Add0~5_sumout ),
	.datac(!\Add0~9_sumout ),
	.datad(!\Add0~13_sumout ),
	.datae(!\LessThan1~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan1~1 .extended_lut = "off";
defparam \LessThan1~1 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \LessThan1~1 .shared_arith = "off";

dffeas fifo_AF(
	.clk(clk_clk),
	.d(\LessThan1~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\fifo_AF~q ),
	.prn(vcc));
defparam fifo_AF.is_wysiwyg = "true";
defparam fifo_AF.power_up = "low";

cyclonev_lcell_comb \fifo_rd~1 (
	.dataa(!A_mem_baddr_2),
	.datab(!av_waitrequest1),
	.datac(!av_waitrequest2),
	.datad(!read_latency_shift_reg),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fifo_rd~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_rd~1 .extended_lut = "off";
defparam \fifo_rd~1 .lut_mask = 64'hEFFFEFFFEFFFEFFF;
defparam \fifo_rd~1 .shared_arith = "off";

cyclonev_lcell_comb \ac~0 (
	.dataa(!\ien_AE~0_combout ),
	.datab(!\first_nios2_system_jtag_uart_alt_jtag_atlantic|t_pause~q ),
	.datac(!\first_nios2_system_jtag_uart_alt_jtag_atlantic|t_ena~q ),
	.datad(!ac1),
	.datae(!A_st_data_10),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac~0 .extended_lut = "off";
defparam \ac~0 .lut_mask = 64'hFFFFBFFFFFFFBFFF;
defparam \ac~0 .shared_arith = "off";

cyclonev_lcell_comb \rvalid~0 (
	.dataa(!b_non_empty),
	.datab(!\fifo_rd~1_combout ),
	.datac(!rvalid1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rvalid~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rvalid~0 .extended_lut = "off";
defparam \rvalid~0 .lut_mask = 64'h4747474747474747;
defparam \rvalid~0 .shared_arith = "off";

cyclonev_lcell_comb \woverflow~0 (
	.dataa(!clr_break_line),
	.datab(!d_write),
	.datac(!A_mem_baddr_2),
	.datad(!av_waitrequest1),
	.datae(!av_waitrequest2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\woverflow~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \woverflow~0 .extended_lut = "off";
defparam \woverflow~0 .lut_mask = 64'hFFF7FFFFFFF7FFFF;
defparam \woverflow~0 .shared_arith = "off";

cyclonev_lcell_comb \woverflow~1 (
	.dataa(!b_full1),
	.datab(!\woverflow~0_combout ),
	.datac(!woverflow1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\woverflow~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \woverflow~1 .extended_lut = "off";
defparam \woverflow~1 .lut_mask = 64'h4747474747474747;
defparam \woverflow~1 .shared_arith = "off";

endmodule

module first_nios2_system_alt_jtag_atlantic (
	r_dat,
	tdo1,
	clr_break_line,
	rst_n,
	t_dav,
	r_val,
	t_pause1,
	rvalid01,
	t_ena1,
	wdata_0,
	wdata_1,
	wdata_2,
	wdata_3,
	wdata_4,
	wdata_5,
	wdata_6,
	wdata_7,
	altera_internal_jtag,
	altera_internal_jtag1,
	state_4,
	splitter_nodes_receive_0_3,
	virtual_ir_scan_reg,
	clr_reg,
	state_3,
	state_8,
	irf_reg_0_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	[7:0] r_dat;
output 	tdo1;
input 	clr_break_line;
input 	rst_n;
input 	t_dav;
input 	r_val;
output 	t_pause1;
output 	rvalid01;
output 	t_ena1;
output 	wdata_0;
output 	wdata_1;
output 	wdata_2;
output 	wdata_3;
output 	wdata_4;
output 	wdata_5;
output 	wdata_6;
output 	wdata_7;
input 	altera_internal_jtag;
input 	altera_internal_jtag1;
input 	state_4;
input 	splitter_nodes_receive_0_3;
input 	virtual_ir_scan_reg;
input 	clr_reg;
input 	state_3;
input 	state_8;
input 	irf_reg_0_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \state~1_combout ;
wire \state~q ;
wire \td_shift[0]~2_combout ;
wire \count[2]~q ;
wire \count[3]~q ;
wire \count[4]~q ;
wire \count[5]~q ;
wire \count[6]~q ;
wire \count[7]~q ;
wire \count[8]~q ;
wire \count[9]~0_combout ;
wire \count[9]~q ;
wire \count[9]~_wirecell_combout ;
wire \count[0]~q ;
wire \count[1]~q ;
wire \state~0_combout ;
wire \user_saw_rvalid~0_combout ;
wire \user_saw_rvalid~q ;
wire \td_shift[10]~q ;
wire \r_ena1~q ;
wire \r_ena~0_combout ;
wire \rdata[7]~q ;
wire \td_shift~3_combout ;
wire \td_shift[9]~q ;
wire \td_shift~0_combout ;
wire \tck_t_dav~0_combout ;
wire \tck_t_dav~q ;
wire \write_stalled~0_combout ;
wire \write_stalled~1_combout ;
wire \write_stalled~q ;
wire \td_shift~4_combout ;
wire \rdata[0]~q ;
wire \rdata[3]~q ;
wire \rdata[6]~q ;
wire \td_shift~12_combout ;
wire \td_shift[8]~q ;
wire \rdata[5]~q ;
wire \td_shift~11_combout ;
wire \td_shift[7]~q ;
wire \rdata[4]~q ;
wire \td_shift~10_combout ;
wire \td_shift[6]~q ;
wire \td_shift~9_combout ;
wire \td_shift[5]~q ;
wire \rdata[2]~q ;
wire \td_shift~8_combout ;
wire \td_shift[4]~q ;
wire \rdata[1]~q ;
wire \td_shift~7_combout ;
wire \td_shift[3]~q ;
wire \td_shift~6_combout ;
wire \td_shift[2]~q ;
wire \td_shift~5_combout ;
wire \td_shift[1]~q ;
wire \read_req~q ;
wire \read~0_combout ;
wire \read~q ;
wire \read1~q ;
wire \read2~q ;
wire \always2~0_combout ;
wire \rst2~q ;
wire \rvalid0~0_combout ;
wire \rvalid0~q ;
wire \rvalid~q ;
wire \td_shift~1_combout ;
wire \td_shift[0]~q ;
wire \jupdate~0_combout ;
wire \jupdate~q ;
wire \jupdate1~q ;
wire \jupdate2~q ;
wire \always2~1_combout ;
wire \write~1_combout ;
wire \write~0_combout ;
wire \write~q ;
wire \write1~q ;
wire \write2~q ;
wire \always2~2_combout ;
wire \write_valid~q ;
wire \t_pause~0_combout ;
wire \t_ena~0_combout ;


dffeas tdo(
	.clk(!altera_internal_jtag),
	.d(\td_shift[0]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(tdo1),
	.prn(vcc));
defparam tdo.is_wysiwyg = "true";
defparam tdo.power_up = "low";

dffeas t_pause(
	.clk(clk),
	.d(\t_pause~0_combout ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(t_pause1),
	.prn(vcc));
defparam t_pause.is_wysiwyg = "true";
defparam t_pause.power_up = "low";

cyclonev_lcell_comb \rvalid0~1 (
	.dataa(!\rvalid0~q ),
	.datab(!\r_ena~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rvalid01),
	.sumout(),
	.cout(),
	.shareout());
defparam \rvalid0~1 .extended_lut = "off";
defparam \rvalid0~1 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \rvalid0~1 .shared_arith = "off";

dffeas t_ena(
	.clk(clk),
	.d(\t_ena~0_combout ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(t_ena1),
	.prn(vcc));
defparam t_ena.is_wysiwyg = "true";
defparam t_ena.power_up = "low";

dffeas \wdata[0] (
	.clk(altera_internal_jtag),
	.d(altera_internal_jtag1),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_stalled~1_combout ),
	.q(wdata_0),
	.prn(vcc));
defparam \wdata[0] .is_wysiwyg = "true";
defparam \wdata[0] .power_up = "low";

dffeas \wdata[1] (
	.clk(altera_internal_jtag),
	.d(\td_shift[5]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write~0_combout ),
	.q(wdata_1),
	.prn(vcc));
defparam \wdata[1] .is_wysiwyg = "true";
defparam \wdata[1] .power_up = "low";

dffeas \wdata[2] (
	.clk(altera_internal_jtag),
	.d(\td_shift[6]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write~0_combout ),
	.q(wdata_2),
	.prn(vcc));
defparam \wdata[2] .is_wysiwyg = "true";
defparam \wdata[2] .power_up = "low";

dffeas \wdata[3] (
	.clk(altera_internal_jtag),
	.d(\td_shift[7]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write~0_combout ),
	.q(wdata_3),
	.prn(vcc));
defparam \wdata[3] .is_wysiwyg = "true";
defparam \wdata[3] .power_up = "low";

dffeas \wdata[4] (
	.clk(altera_internal_jtag),
	.d(\td_shift[8]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write~0_combout ),
	.q(wdata_4),
	.prn(vcc));
defparam \wdata[4] .is_wysiwyg = "true";
defparam \wdata[4] .power_up = "low";

dffeas \wdata[5] (
	.clk(altera_internal_jtag),
	.d(\td_shift[9]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write~0_combout ),
	.q(wdata_5),
	.prn(vcc));
defparam \wdata[5] .is_wysiwyg = "true";
defparam \wdata[5] .power_up = "low";

dffeas \wdata[6] (
	.clk(altera_internal_jtag),
	.d(\td_shift[10]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write~0_combout ),
	.q(wdata_6),
	.prn(vcc));
defparam \wdata[6] .is_wysiwyg = "true";
defparam \wdata[6] .power_up = "low";

dffeas \wdata[7] (
	.clk(altera_internal_jtag),
	.d(altera_internal_jtag1),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write~0_combout ),
	.q(wdata_7),
	.prn(vcc));
defparam \wdata[7] .is_wysiwyg = "true";
defparam \wdata[7] .power_up = "low";

cyclonev_lcell_comb \state~1 (
	.dataa(!virtual_ir_scan_reg),
	.datab(!splitter_nodes_receive_0_3),
	.datac(!state_3),
	.datad(!state_4),
	.datae(!\state~q ),
	.dataf(!altera_internal_jtag1),
	.datag(!irf_reg_0_1),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~1 .extended_lut = "on";
defparam \state~1 .lut_mask = 64'hFF6FFF6FFF6FFF6F;
defparam \state~1 .shared_arith = "off";

dffeas state(
	.clk(altera_internal_jtag),
	.d(\state~1_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state~q ),
	.prn(vcc));
defparam state.is_wysiwyg = "true";
defparam state.power_up = "low";

cyclonev_lcell_comb \td_shift[0]~2 (
	.dataa(!state_4),
	.datab(!splitter_nodes_receive_0_3),
	.datac(!virtual_ir_scan_reg),
	.datad(!state_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\td_shift[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \td_shift[0]~2 .extended_lut = "off";
defparam \td_shift[0]~2 .lut_mask = 64'hF7FFF7FFF7FFF7FF;
defparam \td_shift[0]~2 .shared_arith = "off";

dffeas \count[2] (
	.clk(altera_internal_jtag),
	.d(\count[1]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(!state_4),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\count[2]~q ),
	.prn(vcc));
defparam \count[2] .is_wysiwyg = "true";
defparam \count[2] .power_up = "low";

dffeas \count[3] (
	.clk(altera_internal_jtag),
	.d(\count[2]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(!state_4),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\count[3]~q ),
	.prn(vcc));
defparam \count[3] .is_wysiwyg = "true";
defparam \count[3] .power_up = "low";

dffeas \count[4] (
	.clk(altera_internal_jtag),
	.d(\count[3]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(!state_4),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\count[4]~q ),
	.prn(vcc));
defparam \count[4] .is_wysiwyg = "true";
defparam \count[4] .power_up = "low";

dffeas \count[5] (
	.clk(altera_internal_jtag),
	.d(\count[4]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(!state_4),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\count[5]~q ),
	.prn(vcc));
defparam \count[5] .is_wysiwyg = "true";
defparam \count[5] .power_up = "low";

dffeas \count[6] (
	.clk(altera_internal_jtag),
	.d(\count[5]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(!state_4),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\count[6]~q ),
	.prn(vcc));
defparam \count[6] .is_wysiwyg = "true";
defparam \count[6] .power_up = "low";

dffeas \count[7] (
	.clk(altera_internal_jtag),
	.d(\count[6]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(!state_4),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\count[7]~q ),
	.prn(vcc));
defparam \count[7] .is_wysiwyg = "true";
defparam \count[7] .power_up = "low";

dffeas \count[8] (
	.clk(altera_internal_jtag),
	.d(\count[7]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(!state_4),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\count[8]~q ),
	.prn(vcc));
defparam \count[8] .is_wysiwyg = "true";
defparam \count[8] .power_up = "low";

cyclonev_lcell_comb \count[9]~0 (
	.dataa(!irf_reg_0_1),
	.datab(!\state~q ),
	.datac(!altera_internal_jtag1),
	.datad(!state_4),
	.datae(!\count[8]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\count[9]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \count[9]~0 .extended_lut = "off";
defparam \count[9]~0 .lut_mask = 64'hFFFFFFF7FFFFFFF7;
defparam \count[9]~0 .shared_arith = "off";

dffeas \count[9] (
	.clk(altera_internal_jtag),
	.d(\count[9]~0_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\count[9]~q ),
	.prn(vcc));
defparam \count[9] .is_wysiwyg = "true";
defparam \count[9] .power_up = "low";

cyclonev_lcell_comb \count[9]~_wirecell (
	.dataa(!\count[9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\count[9]~_wirecell_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \count[9]~_wirecell .extended_lut = "off";
defparam \count[9]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \count[9]~_wirecell .shared_arith = "off";

dffeas \count[0] (
	.clk(altera_internal_jtag),
	.d(\count[9]~_wirecell_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(!state_4),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\count[0]~q ),
	.prn(vcc));
defparam \count[0] .is_wysiwyg = "true";
defparam \count[0] .power_up = "low";

dffeas \count[1] (
	.clk(altera_internal_jtag),
	.d(\count[0]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(!state_4),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\count[1]~q ),
	.prn(vcc));
defparam \count[1] .is_wysiwyg = "true";
defparam \count[1] .power_up = "low";

cyclonev_lcell_comb \state~0 (
	.dataa(!state_4),
	.datab(!splitter_nodes_receive_0_3),
	.datac(!virtual_ir_scan_reg),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~0 .extended_lut = "off";
defparam \state~0 .lut_mask = 64'hF7F7F7F7F7F7F7F7;
defparam \state~0 .shared_arith = "off";

cyclonev_lcell_comb \user_saw_rvalid~0 (
	.dataa(!irf_reg_0_1),
	.datab(!\td_shift[0]~q ),
	.datac(!\state~q ),
	.datad(!\user_saw_rvalid~q ),
	.datae(!\state~0_combout ),
	.dataf(!\count[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\user_saw_rvalid~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \user_saw_rvalid~0 .extended_lut = "off";
defparam \user_saw_rvalid~0 .lut_mask = 64'h7BFFB7FFB7FF7BFF;
defparam \user_saw_rvalid~0 .shared_arith = "off";

dffeas user_saw_rvalid(
	.clk(altera_internal_jtag),
	.d(\user_saw_rvalid~0_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\user_saw_rvalid~q ),
	.prn(vcc));
defparam user_saw_rvalid.is_wysiwyg = "true";
defparam user_saw_rvalid.power_up = "low";

dffeas \td_shift[10] (
	.clk(altera_internal_jtag),
	.d(altera_internal_jtag1),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(!state_4),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\td_shift[10]~q ),
	.prn(vcc));
defparam \td_shift[10] .is_wysiwyg = "true";
defparam \td_shift[10] .power_up = "low";

dffeas r_ena1(
	.clk(clk),
	.d(rvalid01),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\r_ena1~q ),
	.prn(vcc));
defparam r_ena1.is_wysiwyg = "true";
defparam r_ena1.power_up = "low";

cyclonev_lcell_comb \r_ena~0 (
	.dataa(!r_val),
	.datab(!\r_ena1~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\r_ena~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \r_ena~0 .extended_lut = "off";
defparam \r_ena~0 .lut_mask = 64'h7777777777777777;
defparam \r_ena~0 .shared_arith = "off";

dffeas \rdata[7] (
	.clk(clk),
	.d(r_dat[7]),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\r_ena~0_combout ),
	.q(\rdata[7]~q ),
	.prn(vcc));
defparam \rdata[7] .is_wysiwyg = "true";
defparam \rdata[7] .power_up = "low";

cyclonev_lcell_comb \td_shift~3 (
	.dataa(!\count[9]~q ),
	.datab(!\td_shift[10]~q ),
	.datac(!\rdata[7]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\td_shift~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \td_shift~3 .extended_lut = "off";
defparam \td_shift~3 .lut_mask = 64'h2727272727272727;
defparam \td_shift~3 .shared_arith = "off";

dffeas \td_shift[9] (
	.clk(altera_internal_jtag),
	.d(\td_shift~3_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(!state_4),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\td_shift[9]~q ),
	.prn(vcc));
defparam \td_shift[9] .is_wysiwyg = "true";
defparam \td_shift[9] .power_up = "low";

cyclonev_lcell_comb \td_shift~0 (
	.dataa(!irf_reg_0_1),
	.datab(!\state~q ),
	.datac(!\count[1]~q ),
	.datad(!\user_saw_rvalid~q ),
	.datae(!\td_shift[9]~q ),
	.dataf(!altera_internal_jtag1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\td_shift~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \td_shift~0 .extended_lut = "off";
defparam \td_shift~0 .lut_mask = 64'hFFFFBF8FFFFFFFFF;
defparam \td_shift~0 .shared_arith = "off";

cyclonev_lcell_comb \tck_t_dav~0 (
	.dataa(!t_dav),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\tck_t_dav~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \tck_t_dav~0 .extended_lut = "off";
defparam \tck_t_dav~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \tck_t_dav~0 .shared_arith = "off";

dffeas tck_t_dav(
	.clk(altera_internal_jtag),
	.d(\tck_t_dav~0_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\tck_t_dav~q ),
	.prn(vcc));
defparam tck_t_dav.is_wysiwyg = "true";
defparam tck_t_dav.power_up = "low";

cyclonev_lcell_comb \write_stalled~0 (
	.dataa(!altera_internal_jtag1),
	.datab(!\tck_t_dav~q ),
	.datac(!\td_shift[10]~q ),
	.datad(!\write_stalled~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\write_stalled~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \write_stalled~0 .extended_lut = "off";
defparam \write_stalled~0 .lut_mask = 64'hEFFFEFFFEFFFEFFF;
defparam \write_stalled~0 .shared_arith = "off";

cyclonev_lcell_comb \write_stalled~1 (
	.dataa(!irf_reg_0_1),
	.datab(!\state~q ),
	.datac(!\count[1]~q ),
	.datad(!state_4),
	.datae(!splitter_nodes_receive_0_3),
	.dataf(!virtual_ir_scan_reg),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\write_stalled~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \write_stalled~1 .extended_lut = "off";
defparam \write_stalled~1 .lut_mask = 64'hFFFFFFFFBFFFFFFF;
defparam \write_stalled~1 .shared_arith = "off";

dffeas write_stalled(
	.clk(altera_internal_jtag),
	.d(\write_stalled~0_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_stalled~1_combout ),
	.q(\write_stalled~q ),
	.prn(vcc));
defparam write_stalled.is_wysiwyg = "true";
defparam write_stalled.power_up = "low";

cyclonev_lcell_comb \td_shift~4 (
	.dataa(!irf_reg_0_1),
	.datab(!\state~q ),
	.datac(!\count[1]~q ),
	.datad(!\user_saw_rvalid~q ),
	.datae(!\td_shift[9]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\td_shift~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \td_shift~4 .extended_lut = "off";
defparam \td_shift~4 .lut_mask = 64'hFFFFFFBFFFFFFFBF;
defparam \td_shift~4 .shared_arith = "off";

dffeas \rdata[0] (
	.clk(clk),
	.d(r_dat[0]),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\r_ena~0_combout ),
	.q(\rdata[0]~q ),
	.prn(vcc));
defparam \rdata[0] .is_wysiwyg = "true";
defparam \rdata[0] .power_up = "low";

dffeas \rdata[3] (
	.clk(clk),
	.d(r_dat[3]),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\r_ena~0_combout ),
	.q(\rdata[3]~q ),
	.prn(vcc));
defparam \rdata[3] .is_wysiwyg = "true";
defparam \rdata[3] .power_up = "low";

dffeas \rdata[6] (
	.clk(clk),
	.d(r_dat[6]),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\r_ena~0_combout ),
	.q(\rdata[6]~q ),
	.prn(vcc));
defparam \rdata[6] .is_wysiwyg = "true";
defparam \rdata[6] .power_up = "low";

cyclonev_lcell_comb \td_shift~12 (
	.dataa(!\td_shift[9]~q ),
	.datab(!\count[9]~q ),
	.datac(!\rdata[6]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\td_shift~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \td_shift~12 .extended_lut = "off";
defparam \td_shift~12 .lut_mask = 64'h4747474747474747;
defparam \td_shift~12 .shared_arith = "off";

dffeas \td_shift[8] (
	.clk(altera_internal_jtag),
	.d(\td_shift~12_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(!state_4),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\td_shift[8]~q ),
	.prn(vcc));
defparam \td_shift[8] .is_wysiwyg = "true";
defparam \td_shift[8] .power_up = "low";

dffeas \rdata[5] (
	.clk(clk),
	.d(r_dat[5]),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\r_ena~0_combout ),
	.q(\rdata[5]~q ),
	.prn(vcc));
defparam \rdata[5] .is_wysiwyg = "true";
defparam \rdata[5] .power_up = "low";

cyclonev_lcell_comb \td_shift~11 (
	.dataa(!\count[9]~q ),
	.datab(!state_4),
	.datac(!\td_shift~4_combout ),
	.datad(!\td_shift[8]~q ),
	.datae(!\rdata[5]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\td_shift~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \td_shift~11 .extended_lut = "off";
defparam \td_shift~11 .lut_mask = 64'hB1FFFFFFB1FFFFFF;
defparam \td_shift~11 .shared_arith = "off";

dffeas \td_shift[7] (
	.clk(altera_internal_jtag),
	.d(\td_shift~11_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\td_shift[7]~q ),
	.prn(vcc));
defparam \td_shift[7] .is_wysiwyg = "true";
defparam \td_shift[7] .power_up = "low";

dffeas \rdata[4] (
	.clk(clk),
	.d(r_dat[4]),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\r_ena~0_combout ),
	.q(\rdata[4]~q ),
	.prn(vcc));
defparam \rdata[4] .is_wysiwyg = "true";
defparam \rdata[4] .power_up = "low";

cyclonev_lcell_comb \td_shift~10 (
	.dataa(!irf_reg_0_1),
	.datab(!\count[9]~q ),
	.datac(!state_4),
	.datad(!\td_shift~4_combout ),
	.datae(!\td_shift[7]~q ),
	.dataf(!\rdata[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\td_shift~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \td_shift~10 .extended_lut = "off";
defparam \td_shift~10 .lut_mask = 64'hFF7DFFFFFFFFFFFF;
defparam \td_shift~10 .shared_arith = "off";

dffeas \td_shift[6] (
	.clk(altera_internal_jtag),
	.d(\td_shift~10_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\td_shift[6]~q ),
	.prn(vcc));
defparam \td_shift[6] .is_wysiwyg = "true";
defparam \td_shift[6] .power_up = "low";

cyclonev_lcell_comb \td_shift~9 (
	.dataa(!irf_reg_0_1),
	.datab(!\count[9]~q ),
	.datac(!state_4),
	.datad(!\td_shift~4_combout ),
	.datae(!\rdata[3]~q ),
	.dataf(!\td_shift[6]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\td_shift~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \td_shift~9 .extended_lut = "off";
defparam \td_shift~9 .lut_mask = 64'hFF7DFFFFFFFFFFFF;
defparam \td_shift~9 .shared_arith = "off";

dffeas \td_shift[5] (
	.clk(altera_internal_jtag),
	.d(\td_shift~9_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\td_shift[5]~q ),
	.prn(vcc));
defparam \td_shift[5] .is_wysiwyg = "true";
defparam \td_shift[5] .power_up = "low";

dffeas \rdata[2] (
	.clk(clk),
	.d(r_dat[2]),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\r_ena~0_combout ),
	.q(\rdata[2]~q ),
	.prn(vcc));
defparam \rdata[2] .is_wysiwyg = "true";
defparam \rdata[2] .power_up = "low";

cyclonev_lcell_comb \td_shift~8 (
	.dataa(!\count[9]~q ),
	.datab(!state_4),
	.datac(!\td_shift~4_combout ),
	.datad(!\td_shift[5]~q ),
	.datae(!\rdata[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\td_shift~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \td_shift~8 .extended_lut = "off";
defparam \td_shift~8 .lut_mask = 64'hB1FFFFFFB1FFFFFF;
defparam \td_shift~8 .shared_arith = "off";

dffeas \td_shift[4] (
	.clk(altera_internal_jtag),
	.d(\td_shift~8_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\td_shift[4]~q ),
	.prn(vcc));
defparam \td_shift[4] .is_wysiwyg = "true";
defparam \td_shift[4] .power_up = "low";

dffeas \rdata[1] (
	.clk(clk),
	.d(r_dat[1]),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\r_ena~0_combout ),
	.q(\rdata[1]~q ),
	.prn(vcc));
defparam \rdata[1] .is_wysiwyg = "true";
defparam \rdata[1] .power_up = "low";

cyclonev_lcell_comb \td_shift~7 (
	.dataa(!\count[9]~q ),
	.datab(!state_4),
	.datac(!\td_shift~4_combout ),
	.datad(!\td_shift[4]~q ),
	.datae(!\rdata[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\td_shift~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \td_shift~7 .extended_lut = "off";
defparam \td_shift~7 .lut_mask = 64'hB1FFFFFFB1FFFFFF;
defparam \td_shift~7 .shared_arith = "off";

dffeas \td_shift[3] (
	.clk(altera_internal_jtag),
	.d(\td_shift~7_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\td_shift[3]~q ),
	.prn(vcc));
defparam \td_shift[3] .is_wysiwyg = "true";
defparam \td_shift[3] .power_up = "low";

cyclonev_lcell_comb \td_shift~6 (
	.dataa(!irf_reg_0_1),
	.datab(!\count[9]~q ),
	.datac(!state_4),
	.datad(!\td_shift~4_combout ),
	.datae(!\rdata[0]~q ),
	.dataf(!\td_shift[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\td_shift~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \td_shift~6 .extended_lut = "off";
defparam \td_shift~6 .lut_mask = 64'hFF7DFFFFFFFFFFFF;
defparam \td_shift~6 .shared_arith = "off";

dffeas \td_shift[2] (
	.clk(altera_internal_jtag),
	.d(\td_shift~6_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\td_shift[2]~q ),
	.prn(vcc));
defparam \td_shift[2] .is_wysiwyg = "true";
defparam \td_shift[2] .power_up = "low";

cyclonev_lcell_comb \td_shift~5 (
	.dataa(!irf_reg_0_1),
	.datab(!\count[9]~q ),
	.datac(!state_4),
	.datad(!\write_stalled~q ),
	.datae(!\td_shift~4_combout ),
	.dataf(!\td_shift[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\td_shift~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \td_shift~5 .extended_lut = "off";
defparam \td_shift~5 .lut_mask = 64'hFFFF7DFFFFFFFFFF;
defparam \td_shift~5 .shared_arith = "off";

dffeas \td_shift[1] (
	.clk(altera_internal_jtag),
	.d(\td_shift~5_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\td_shift[1]~q ),
	.prn(vcc));
defparam \td_shift[1] .is_wysiwyg = "true";
defparam \td_shift[1] .power_up = "low";

dffeas read_req(
	.clk(altera_internal_jtag),
	.d(\td_shift[9]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_stalled~1_combout ),
	.q(\read_req~q ),
	.prn(vcc));
defparam read_req.is_wysiwyg = "true";
defparam read_req.power_up = "low";

cyclonev_lcell_comb \read~0 (
	.dataa(!\read~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read~0 .extended_lut = "off";
defparam \read~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \read~0 .shared_arith = "off";

dffeas read(
	.clk(altera_internal_jtag),
	.d(\read~0_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_stalled~1_combout ),
	.q(\read~q ),
	.prn(vcc));
defparam read.is_wysiwyg = "true";
defparam read.power_up = "low";

dffeas read1(
	.clk(clk),
	.d(\read~q ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\read1~q ),
	.prn(vcc));
defparam read1.is_wysiwyg = "true";
defparam read1.power_up = "low";

dffeas read2(
	.clk(clk),
	.d(\read1~q ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\read2~q ),
	.prn(vcc));
defparam read2.is_wysiwyg = "true";
defparam read2.power_up = "low";

cyclonev_lcell_comb \always2~0 (
	.dataa(!\read1~q ),
	.datab(!\read2~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always2~0 .extended_lut = "off";
defparam \always2~0 .lut_mask = 64'h6666666666666666;
defparam \always2~0 .shared_arith = "off";

dffeas rst2(
	.clk(clk),
	.d(clr_break_line),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rst2~q ),
	.prn(vcc));
defparam rst2.is_wysiwyg = "true";
defparam rst2.power_up = "low";

cyclonev_lcell_comb \rvalid0~0 (
	.dataa(!\user_saw_rvalid~q ),
	.datab(!\rvalid0~q ),
	.datac(!\r_ena~0_combout ),
	.datad(!\read_req~q ),
	.datae(!\always2~0_combout ),
	.dataf(!\rst2~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rvalid0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rvalid0~0 .extended_lut = "off";
defparam \rvalid0~0 .lut_mask = 64'hFFFFFFFFFFFFFFBF;
defparam \rvalid0~0 .shared_arith = "off";

dffeas rvalid0(
	.clk(clk),
	.d(\rvalid0~0_combout ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rvalid0~q ),
	.prn(vcc));
defparam rvalid0.is_wysiwyg = "true";
defparam rvalid0.power_up = "low";

dffeas rvalid(
	.clk(clk),
	.d(\rvalid0~q ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rvalid~q ),
	.prn(vcc));
defparam rvalid.is_wysiwyg = "true";
defparam rvalid.power_up = "low";

cyclonev_lcell_comb \td_shift~1 (
	.dataa(!\state~q ),
	.datab(!\td_shift~0_combout ),
	.datac(!\tck_t_dav~q ),
	.datad(!\td_shift[1]~q ),
	.datae(!\count[9]~q ),
	.dataf(!\rvalid~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\td_shift~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \td_shift~1 .extended_lut = "off";
defparam \td_shift~1 .lut_mask = 64'hBFFFEFFFFFFFFFFF;
defparam \td_shift~1 .shared_arith = "off";

dffeas \td_shift[0] (
	.clk(altera_internal_jtag),
	.d(\td_shift~1_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(!state_4),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\td_shift[0]~q ),
	.prn(vcc));
defparam \td_shift[0] .is_wysiwyg = "true";
defparam \td_shift[0] .power_up = "low";

cyclonev_lcell_comb \jupdate~0 (
	.dataa(!irf_reg_0_1),
	.datab(!splitter_nodes_receive_0_3),
	.datac(!virtual_ir_scan_reg),
	.datad(!\jupdate~q ),
	.datae(!state_8),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\jupdate~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \jupdate~0 .extended_lut = "off";
defparam \jupdate~0 .lut_mask = 64'h9669699696696996;
defparam \jupdate~0 .shared_arith = "off";

dffeas jupdate(
	.clk(!altera_internal_jtag),
	.d(\jupdate~0_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jupdate~q ),
	.prn(vcc));
defparam jupdate.is_wysiwyg = "true";
defparam jupdate.power_up = "low";

dffeas jupdate1(
	.clk(clk),
	.d(\jupdate~q ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jupdate1~q ),
	.prn(vcc));
defparam jupdate1.is_wysiwyg = "true";
defparam jupdate1.power_up = "low";

dffeas jupdate2(
	.clk(clk),
	.d(\jupdate1~q ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jupdate2~q ),
	.prn(vcc));
defparam jupdate2.is_wysiwyg = "true";
defparam jupdate2.power_up = "low";

cyclonev_lcell_comb \always2~1 (
	.dataa(!\jupdate1~q ),
	.datab(!\jupdate2~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always2~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always2~1 .extended_lut = "off";
defparam \always2~1 .lut_mask = 64'h6666666666666666;
defparam \always2~1 .shared_arith = "off";

cyclonev_lcell_comb \write~1 (
	.dataa(!\write~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\write~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \write~1 .extended_lut = "off";
defparam \write~1 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \write~1 .shared_arith = "off";

cyclonev_lcell_comb \write~0 (
	.dataa(!irf_reg_0_1),
	.datab(!\state~q ),
	.datac(!state_4),
	.datad(!splitter_nodes_receive_0_3),
	.datae(!virtual_ir_scan_reg),
	.dataf(!\count[8]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\write~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \write~0 .extended_lut = "off";
defparam \write~0 .lut_mask = 64'hFFFFBFFFFFFFFFFF;
defparam \write~0 .shared_arith = "off";

dffeas write(
	.clk(altera_internal_jtag),
	.d(\write~1_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write~0_combout ),
	.q(\write~q ),
	.prn(vcc));
defparam write.is_wysiwyg = "true";
defparam write.power_up = "low";

dffeas write1(
	.clk(clk),
	.d(\write~q ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\write1~q ),
	.prn(vcc));
defparam write1.is_wysiwyg = "true";
defparam write1.power_up = "low";

dffeas write2(
	.clk(clk),
	.d(\write1~q ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\write2~q ),
	.prn(vcc));
defparam write2.is_wysiwyg = "true";
defparam write2.power_up = "low";

cyclonev_lcell_comb \always2~2 (
	.dataa(!\write1~q ),
	.datab(!\write2~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always2~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always2~2 .extended_lut = "off";
defparam \always2~2 .lut_mask = 64'h6666666666666666;
defparam \always2~2 .shared_arith = "off";

dffeas write_valid(
	.clk(altera_internal_jtag),
	.d(\td_shift[10]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_stalled~1_combout ),
	.q(\write_valid~q ),
	.prn(vcc));
defparam write_valid.is_wysiwyg = "true";
defparam write_valid.power_up = "low";

cyclonev_lcell_comb \t_pause~0 (
	.dataa(!t_dav),
	.datab(!\write_stalled~q ),
	.datac(!\rst2~q ),
	.datad(!\always2~1_combout ),
	.datae(!\always2~2_combout ),
	.dataf(!\write_valid~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\t_pause~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \t_pause~0 .extended_lut = "off";
defparam \t_pause~0 .lut_mask = 64'hFFFFFFFF7FFFFFFF;
defparam \t_pause~0 .shared_arith = "off";

cyclonev_lcell_comb \t_ena~0 (
	.dataa(!t_dav),
	.datab(!\write_stalled~q ),
	.datac(!\rst2~q ),
	.datad(!t_ena1),
	.datae(!\always2~2_combout ),
	.dataf(!\write_valid~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\t_ena~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \t_ena~0 .extended_lut = "off";
defparam \t_ena~0 .lut_mask = 64'hEFFFFFFFFFFFFFFF;
defparam \t_ena~0 .shared_arith = "off";

endmodule

module first_nios2_system_first_nios2_system_jtag_uart_scfifo_r (
	q_b_0,
	q_b_1,
	q_b_2,
	q_b_3,
	q_b_4,
	q_b_5,
	q_b_6,
	q_b_7,
	A_mem_baddr_2,
	r_sync_rst,
	read_latency_shift_reg,
	av_waitrequest,
	av_waitrequest1,
	b_full,
	b_non_empty,
	counter_reg_bit_0,
	counter_reg_bit_1,
	fifo_rd,
	t_ena,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_5,
	wr_rfifo,
	wdata_0,
	wdata_1,
	wdata_2,
	wdata_3,
	wdata_4,
	wdata_5,
	wdata_6,
	wdata_7,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_0;
output 	q_b_1;
output 	q_b_2;
output 	q_b_3;
output 	q_b_4;
output 	q_b_5;
output 	q_b_6;
output 	q_b_7;
input 	A_mem_baddr_2;
input 	r_sync_rst;
input 	read_latency_shift_reg;
input 	av_waitrequest;
input 	av_waitrequest1;
output 	b_full;
output 	b_non_empty;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
input 	fifo_rd;
input 	t_ena;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_5;
input 	wr_rfifo;
input 	wdata_0;
input 	wdata_1;
input 	wdata_2;
input 	wdata_3;
input 	wdata_4;
input 	wdata_5;
input 	wdata_6;
input 	wdata_7;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



first_nios2_system_scfifo_1 rfifo(
	.q({q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.A_mem_baddr_2(A_mem_baddr_2),
	.r_sync_rst(r_sync_rst),
	.read_latency_shift_reg(read_latency_shift_reg),
	.av_waitrequest(av_waitrequest),
	.av_waitrequest1(av_waitrequest1),
	.b_full(b_full),
	.b_non_empty(b_non_empty),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_1(counter_reg_bit_1),
	.fifo_rd(fifo_rd),
	.t_ena(t_ena),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_5(counter_reg_bit_5),
	.wrreq(wr_rfifo),
	.data({wdata_7,wdata_6,wdata_5,wdata_4,wdata_3,wdata_2,wdata_1,wdata_0}),
	.clock(clk_clk));

endmodule

module first_nios2_system_scfifo_1 (
	q,
	A_mem_baddr_2,
	r_sync_rst,
	read_latency_shift_reg,
	av_waitrequest,
	av_waitrequest1,
	b_full,
	b_non_empty,
	counter_reg_bit_0,
	counter_reg_bit_1,
	fifo_rd,
	t_ena,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_5,
	wrreq,
	data,
	clock)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q;
input 	A_mem_baddr_2;
input 	r_sync_rst;
input 	read_latency_shift_reg;
input 	av_waitrequest;
input 	av_waitrequest1;
output 	b_full;
output 	b_non_empty;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
input 	fifo_rd;
input 	t_ena;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_5;
input 	wrreq;
input 	[7:0] data;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



first_nios2_system_scfifo_3291 auto_generated(
	.q({q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.A_mem_baddr_2(A_mem_baddr_2),
	.r_sync_rst(r_sync_rst),
	.read_latency_shift_reg(read_latency_shift_reg),
	.av_waitrequest(av_waitrequest),
	.av_waitrequest1(av_waitrequest1),
	.b_full(b_full),
	.b_non_empty(b_non_empty),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_1(counter_reg_bit_1),
	.fifo_rd(fifo_rd),
	.t_ena(t_ena),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_5(counter_reg_bit_5),
	.wrreq(wrreq),
	.data({data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.clock(clock));

endmodule

module first_nios2_system_scfifo_3291 (
	q,
	A_mem_baddr_2,
	r_sync_rst,
	read_latency_shift_reg,
	av_waitrequest,
	av_waitrequest1,
	b_full,
	b_non_empty,
	counter_reg_bit_0,
	counter_reg_bit_1,
	fifo_rd,
	t_ena,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_5,
	wrreq,
	data,
	clock)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q;
input 	A_mem_baddr_2;
input 	r_sync_rst;
input 	read_latency_shift_reg;
input 	av_waitrequest;
input 	av_waitrequest1;
output 	b_full;
output 	b_non_empty;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
input 	fifo_rd;
input 	t_ena;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_5;
input 	wrreq;
input 	[7:0] data;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



first_nios2_system_a_dpfifo_5771 dpfifo(
	.q({q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.A_mem_baddr_2(A_mem_baddr_2),
	.r_sync_rst(r_sync_rst),
	.read_latency_shift_reg(read_latency_shift_reg),
	.av_waitrequest(av_waitrequest),
	.av_waitrequest1(av_waitrequest1),
	.b_full(b_full),
	.b_non_empty(b_non_empty),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_1(counter_reg_bit_1),
	.fifo_rd(fifo_rd),
	.t_ena(t_ena),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_5(counter_reg_bit_5),
	.wreq(wrreq),
	.data({data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.clock(clock));

endmodule

module first_nios2_system_a_dpfifo_5771 (
	q,
	A_mem_baddr_2,
	r_sync_rst,
	read_latency_shift_reg,
	av_waitrequest,
	av_waitrequest1,
	b_full,
	b_non_empty,
	counter_reg_bit_0,
	counter_reg_bit_1,
	fifo_rd,
	t_ena,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_5,
	wreq,
	data,
	clock)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q;
input 	A_mem_baddr_2;
input 	r_sync_rst;
input 	read_latency_shift_reg;
input 	av_waitrequest;
input 	av_waitrequest1;
output 	b_full;
output 	b_non_empty;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
input 	fifo_rd;
input 	t_ena;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_5;
input 	wreq;
input 	[7:0] data;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wr_ptr|counter_reg_bit[0]~q ;
wire \wr_ptr|counter_reg_bit[1]~q ;
wire \wr_ptr|counter_reg_bit[2]~q ;
wire \wr_ptr|counter_reg_bit[3]~q ;
wire \wr_ptr|counter_reg_bit[4]~q ;
wire \wr_ptr|counter_reg_bit[5]~q ;
wire \rd_ptr_count|counter_reg_bit[0]~q ;
wire \rd_ptr_count|counter_reg_bit[1]~q ;
wire \rd_ptr_count|counter_reg_bit[2]~q ;
wire \rd_ptr_count|counter_reg_bit[3]~q ;
wire \rd_ptr_count|counter_reg_bit[4]~q ;
wire \rd_ptr_count|counter_reg_bit[5]~q ;


first_nios2_system_cntr_jgb_1 wr_ptr(
	.r_sync_rst(r_sync_rst),
	.wr_rfifo(wreq),
	.counter_reg_bit_0(\wr_ptr|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\wr_ptr|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\wr_ptr|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\wr_ptr|counter_reg_bit[3]~q ),
	.counter_reg_bit_4(\wr_ptr|counter_reg_bit[4]~q ),
	.counter_reg_bit_5(\wr_ptr|counter_reg_bit[5]~q ),
	.clock(clock));

first_nios2_system_cntr_jgb rd_ptr_count(
	.r_sync_rst(r_sync_rst),
	.fifo_rd(fifo_rd),
	.counter_reg_bit_0(\rd_ptr_count|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\rd_ptr_count|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\rd_ptr_count|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\rd_ptr_count|counter_reg_bit[3]~q ),
	.counter_reg_bit_4(\rd_ptr_count|counter_reg_bit[4]~q ),
	.counter_reg_bit_5(\rd_ptr_count|counter_reg_bit[5]~q ),
	.clock(clock));

first_nios2_system_altsyncram_7pu1 FIFOram(
	.q_b({q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.clocken1(fifo_rd),
	.wren_a(wreq),
	.data_a({data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.address_a({\wr_ptr|counter_reg_bit[5]~q ,\wr_ptr|counter_reg_bit[4]~q ,\wr_ptr|counter_reg_bit[3]~q ,\wr_ptr|counter_reg_bit[2]~q ,\wr_ptr|counter_reg_bit[1]~q ,\wr_ptr|counter_reg_bit[0]~q }),
	.address_b({\rd_ptr_count|counter_reg_bit[5]~q ,\rd_ptr_count|counter_reg_bit[4]~q ,\rd_ptr_count|counter_reg_bit[3]~q ,\rd_ptr_count|counter_reg_bit[2]~q ,\rd_ptr_count|counter_reg_bit[1]~q ,\rd_ptr_count|counter_reg_bit[0]~q }),
	.clock1(clock),
	.clock0(clock));

first_nios2_system_a_fefifo_7cf fifo_state(
	.A_mem_baddr_2(A_mem_baddr_2),
	.r_sync_rst(r_sync_rst),
	.read_latency_shift_reg(read_latency_shift_reg),
	.av_waitrequest(av_waitrequest),
	.av_waitrequest1(av_waitrequest1),
	.b_full1(b_full),
	.b_non_empty1(b_non_empty),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_1(counter_reg_bit_1),
	.fifo_rd(fifo_rd),
	.t_ena(t_ena),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_5(counter_reg_bit_5),
	.wr_rfifo(wreq),
	.clock(clock));

endmodule

module first_nios2_system_a_fefifo_7cf (
	A_mem_baddr_2,
	r_sync_rst,
	read_latency_shift_reg,
	av_waitrequest,
	av_waitrequest1,
	b_full1,
	b_non_empty1,
	counter_reg_bit_0,
	counter_reg_bit_1,
	fifo_rd,
	t_ena,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_5,
	wr_rfifo,
	clock)/* synthesis synthesis_greybox=1 */;
input 	A_mem_baddr_2;
input 	r_sync_rst;
input 	read_latency_shift_reg;
input 	av_waitrequest;
input 	av_waitrequest1;
output 	b_full1;
output 	b_non_empty1;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
input 	fifo_rd;
input 	t_ena;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_5;
input 	wr_rfifo;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \_~2_combout ;
wire \b_full~0_combout ;
wire \b_full~1_combout ;
wire \_~0_combout ;
wire \_~1_combout ;
wire \b_non_empty~0_combout ;


first_nios2_system_cntr_vg7 count_usedw(
	.r_sync_rst(r_sync_rst),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_5(counter_reg_bit_5),
	.wr_rfifo(wr_rfifo),
	._(\_~2_combout ),
	.clock(clock));

cyclonev_lcell_comb \_~2 (
	.dataa(!A_mem_baddr_2),
	.datab(!av_waitrequest),
	.datac(!av_waitrequest1),
	.datad(!read_latency_shift_reg),
	.datae(!b_non_empty1),
	.dataf(!wr_rfifo),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\_~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \_~2 .extended_lut = "off";
defparam \_~2 .lut_mask = 64'h6996966996696996;
defparam \_~2 .shared_arith = "off";

dffeas b_full(
	.clk(clock),
	.d(\b_full~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(b_full1),
	.prn(vcc));
defparam b_full.is_wysiwyg = "true";
defparam b_full.power_up = "low";

dffeas b_non_empty(
	.clk(clock),
	.d(\b_non_empty~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(b_non_empty1),
	.prn(vcc));
defparam b_non_empty.is_wysiwyg = "true";
defparam b_non_empty.power_up = "low";

cyclonev_lcell_comb \b_full~0 (
	.dataa(!b_non_empty1),
	.datab(!counter_reg_bit_4),
	.datac(!counter_reg_bit_3),
	.datad(!counter_reg_bit_2),
	.datae(!counter_reg_bit_5),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\b_full~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \b_full~0 .extended_lut = "off";
defparam \b_full~0 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \b_full~0 .shared_arith = "off";

cyclonev_lcell_comb \b_full~1 (
	.dataa(!b_full1),
	.datab(!counter_reg_bit_0),
	.datac(!counter_reg_bit_1),
	.datad(!fifo_rd),
	.datae(!t_ena),
	.dataf(!\b_full~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\b_full~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \b_full~1 .extended_lut = "off";
defparam \b_full~1 .lut_mask = 64'hFF7FFFFFFFFFFFFF;
defparam \b_full~1 .shared_arith = "off";

cyclonev_lcell_comb \_~0 (
	.dataa(!counter_reg_bit_4),
	.datab(!counter_reg_bit_3),
	.datac(!counter_reg_bit_5),
	.datad(!wr_rfifo),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\_~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \_~0 .extended_lut = "off";
defparam \_~0 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \_~0 .shared_arith = "off";

cyclonev_lcell_comb \_~1 (
	.dataa(!counter_reg_bit_2),
	.datab(!counter_reg_bit_0),
	.datac(!counter_reg_bit_1),
	.datad(!\_~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\_~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \_~1 .extended_lut = "off";
defparam \_~1 .lut_mask = 64'hFBFFFBFFFBFFFBFF;
defparam \_~1 .shared_arith = "off";

cyclonev_lcell_comb \b_non_empty~0 (
	.dataa(!b_full1),
	.datab(!b_non_empty1),
	.datac(!fifo_rd),
	.datad(!t_ena),
	.datae(!\_~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\b_non_empty~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \b_non_empty~0 .extended_lut = "off";
defparam \b_non_empty~0 .lut_mask = 64'hF7FFD5FFF7FFD5FF;
defparam \b_non_empty~0 .shared_arith = "off";

endmodule

module first_nios2_system_cntr_vg7 (
	r_sync_rst,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_5,
	wr_rfifo,
	_,
	clock)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_5;
input 	wr_rfifo;
input 	_;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~sumout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~sumout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~sumout ;
wire \counter_comb_bita3~sumout ;
wire \counter_comb_bita2~sumout ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~sumout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

cyclonev_lcell_comb counter_comb_bita0(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita0~sumout ),
	.cout(\counter_comb_bita0~COUT ),
	.shareout());
defparam counter_comb_bita0.extended_lut = "off";
defparam counter_comb_bita0.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita0.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita1(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_1),
	.datae(gnd),
	.dataf(!wr_rfifo),
	.datag(gnd),
	.cin(\counter_comb_bita0~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita1~sumout ),
	.cout(\counter_comb_bita1~COUT ),
	.shareout());
defparam counter_comb_bita1.extended_lut = "off";
defparam counter_comb_bita1.lut_mask = 64'h000000FF000000FF;
defparam counter_comb_bita1.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita2(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_2),
	.datae(gnd),
	.dataf(!wr_rfifo),
	.datag(gnd),
	.cin(\counter_comb_bita1~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita2~sumout ),
	.cout(\counter_comb_bita2~COUT ),
	.shareout());
defparam counter_comb_bita2.extended_lut = "off";
defparam counter_comb_bita2.lut_mask = 64'h000000FF000000FF;
defparam counter_comb_bita2.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita3(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_3),
	.datae(gnd),
	.dataf(!wr_rfifo),
	.datag(gnd),
	.cin(\counter_comb_bita2~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita3~sumout ),
	.cout(\counter_comb_bita3~COUT ),
	.shareout());
defparam counter_comb_bita3.extended_lut = "off";
defparam counter_comb_bita3.lut_mask = 64'h000000FF000000FF;
defparam counter_comb_bita3.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita4(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_4),
	.datae(gnd),
	.dataf(!wr_rfifo),
	.datag(gnd),
	.cin(\counter_comb_bita3~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita4~sumout ),
	.cout(\counter_comb_bita4~COUT ),
	.shareout());
defparam counter_comb_bita4.extended_lut = "off";
defparam counter_comb_bita4.lut_mask = 64'h000000FF000000FF;
defparam counter_comb_bita4.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita5(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_5),
	.datae(gnd),
	.dataf(!wr_rfifo),
	.datag(gnd),
	.cin(\counter_comb_bita4~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita5~sumout ),
	.cout(),
	.shareout());
defparam counter_comb_bita5.extended_lut = "off";
defparam counter_comb_bita5.lut_mask = 64'h000000FF000000FF;
defparam counter_comb_bita5.shared_arith = "off";

endmodule

module first_nios2_system_altsyncram_7pu1 (
	q_b,
	clocken1,
	wren_a,
	data_a,
	address_a,
	address_b,
	clock1,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q_b;
input 	clocken1;
input 	wren_a;
input 	[7:0] data_a;
input 	[5:0] address_a;
input 	[5:0] address_b;
input 	clock1;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

cyclonev_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk1_core_clock_enable = "ena1";
defparam ram_block1a0.clk1_input_clock_enable = "ena1";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "first_nios2_system_jtag_uart:jtag_uart|first_nios2_system_jtag_uart_scfifo_r:the_first_nios2_system_jtag_uart_scfifo_r|scfifo:rfifo|scfifo_3291:auto_generated|a_dpfifo_5771:dpfifo|altsyncram_7pu1:FIFOram|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 6;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 63;
defparam ram_block1a0.port_a_logical_ram_depth = 64;
defparam ram_block1a0.port_a_logical_ram_width = 8;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock1";
defparam ram_block1a0.port_b_address_width = 6;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "none";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 63;
defparam ram_block1a0.port_b_logical_ram_depth = 64;
defparam ram_block1a0.port_b_logical_ram_width = 8;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock1";
defparam ram_block1a0.ram_block_type = "auto";

cyclonev_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk1_core_clock_enable = "ena1";
defparam ram_block1a1.clk1_input_clock_enable = "ena1";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "first_nios2_system_jtag_uart:jtag_uart|first_nios2_system_jtag_uart_scfifo_r:the_first_nios2_system_jtag_uart_scfifo_r|scfifo:rfifo|scfifo_3291:auto_generated|a_dpfifo_5771:dpfifo|altsyncram_7pu1:FIFOram|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 6;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 63;
defparam ram_block1a1.port_a_logical_ram_depth = 64;
defparam ram_block1a1.port_a_logical_ram_width = 8;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock1";
defparam ram_block1a1.port_b_address_width = 6;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "none";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 63;
defparam ram_block1a1.port_b_logical_ram_depth = 64;
defparam ram_block1a1.port_b_logical_ram_width = 8;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock1";
defparam ram_block1a1.ram_block_type = "auto";

cyclonev_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk1_core_clock_enable = "ena1";
defparam ram_block1a2.clk1_input_clock_enable = "ena1";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "first_nios2_system_jtag_uart:jtag_uart|first_nios2_system_jtag_uart_scfifo_r:the_first_nios2_system_jtag_uart_scfifo_r|scfifo:rfifo|scfifo_3291:auto_generated|a_dpfifo_5771:dpfifo|altsyncram_7pu1:FIFOram|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 6;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 63;
defparam ram_block1a2.port_a_logical_ram_depth = 64;
defparam ram_block1a2.port_a_logical_ram_width = 8;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock1";
defparam ram_block1a2.port_b_address_width = 6;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "none";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 63;
defparam ram_block1a2.port_b_logical_ram_depth = 64;
defparam ram_block1a2.port_b_logical_ram_width = 8;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock1";
defparam ram_block1a2.ram_block_type = "auto";

cyclonev_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk1_core_clock_enable = "ena1";
defparam ram_block1a3.clk1_input_clock_enable = "ena1";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "first_nios2_system_jtag_uart:jtag_uart|first_nios2_system_jtag_uart_scfifo_r:the_first_nios2_system_jtag_uart_scfifo_r|scfifo:rfifo|scfifo_3291:auto_generated|a_dpfifo_5771:dpfifo|altsyncram_7pu1:FIFOram|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 6;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 63;
defparam ram_block1a3.port_a_logical_ram_depth = 64;
defparam ram_block1a3.port_a_logical_ram_width = 8;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock1";
defparam ram_block1a3.port_b_address_width = 6;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "none";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 63;
defparam ram_block1a3.port_b_logical_ram_depth = 64;
defparam ram_block1a3.port_b_logical_ram_width = 8;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock1";
defparam ram_block1a3.ram_block_type = "auto";

cyclonev_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk1_core_clock_enable = "ena1";
defparam ram_block1a4.clk1_input_clock_enable = "ena1";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "first_nios2_system_jtag_uart:jtag_uart|first_nios2_system_jtag_uart_scfifo_r:the_first_nios2_system_jtag_uart_scfifo_r|scfifo:rfifo|scfifo_3291:auto_generated|a_dpfifo_5771:dpfifo|altsyncram_7pu1:FIFOram|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 6;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 63;
defparam ram_block1a4.port_a_logical_ram_depth = 64;
defparam ram_block1a4.port_a_logical_ram_width = 8;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock1";
defparam ram_block1a4.port_b_address_width = 6;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "none";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 63;
defparam ram_block1a4.port_b_logical_ram_depth = 64;
defparam ram_block1a4.port_b_logical_ram_width = 8;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock1";
defparam ram_block1a4.ram_block_type = "auto";

cyclonev_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk1_core_clock_enable = "ena1";
defparam ram_block1a5.clk1_input_clock_enable = "ena1";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "first_nios2_system_jtag_uart:jtag_uart|first_nios2_system_jtag_uart_scfifo_r:the_first_nios2_system_jtag_uart_scfifo_r|scfifo:rfifo|scfifo_3291:auto_generated|a_dpfifo_5771:dpfifo|altsyncram_7pu1:FIFOram|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 6;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 63;
defparam ram_block1a5.port_a_logical_ram_depth = 64;
defparam ram_block1a5.port_a_logical_ram_width = 8;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 6;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "none";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 63;
defparam ram_block1a5.port_b_logical_ram_depth = 64;
defparam ram_block1a5.port_b_logical_ram_width = 8;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";

cyclonev_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk1_core_clock_enable = "ena1";
defparam ram_block1a6.clk1_input_clock_enable = "ena1";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "first_nios2_system_jtag_uart:jtag_uart|first_nios2_system_jtag_uart_scfifo_r:the_first_nios2_system_jtag_uart_scfifo_r|scfifo:rfifo|scfifo_3291:auto_generated|a_dpfifo_5771:dpfifo|altsyncram_7pu1:FIFOram|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 6;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 63;
defparam ram_block1a6.port_a_logical_ram_depth = 64;
defparam ram_block1a6.port_a_logical_ram_width = 8;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 6;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "none";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 63;
defparam ram_block1a6.port_b_logical_ram_depth = 64;
defparam ram_block1a6.port_b_logical_ram_width = 8;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";

cyclonev_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk1_core_clock_enable = "ena1";
defparam ram_block1a7.clk1_input_clock_enable = "ena1";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "first_nios2_system_jtag_uart:jtag_uart|first_nios2_system_jtag_uart_scfifo_r:the_first_nios2_system_jtag_uart_scfifo_r|scfifo:rfifo|scfifo_3291:auto_generated|a_dpfifo_5771:dpfifo|altsyncram_7pu1:FIFOram|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 6;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 63;
defparam ram_block1a7.port_a_logical_ram_depth = 64;
defparam ram_block1a7.port_a_logical_ram_width = 8;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 6;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "none";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 63;
defparam ram_block1a7.port_b_logical_ram_depth = 64;
defparam ram_block1a7.port_b_logical_ram_width = 8;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";

endmodule

module first_nios2_system_cntr_jgb (
	r_sync_rst,
	fifo_rd,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	counter_reg_bit_5,
	clock)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
input 	fifo_rd;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
output 	counter_reg_bit_5;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~sumout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~sumout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~sumout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~sumout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~sumout ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~sumout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_rd),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_rd),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_rd),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_rd),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_rd),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_rd),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

cyclonev_lcell_comb counter_comb_bita0(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita0~sumout ),
	.cout(\counter_comb_bita0~COUT ),
	.shareout());
defparam counter_comb_bita0.extended_lut = "off";
defparam counter_comb_bita0.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita0.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita1(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita0~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita1~sumout ),
	.cout(\counter_comb_bita1~COUT ),
	.shareout());
defparam counter_comb_bita1.extended_lut = "off";
defparam counter_comb_bita1.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita1.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita2(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita1~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita2~sumout ),
	.cout(\counter_comb_bita2~COUT ),
	.shareout());
defparam counter_comb_bita2.extended_lut = "off";
defparam counter_comb_bita2.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita2.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita3(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita2~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita3~sumout ),
	.cout(\counter_comb_bita3~COUT ),
	.shareout());
defparam counter_comb_bita3.extended_lut = "off";
defparam counter_comb_bita3.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita3.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita4(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita3~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita4~sumout ),
	.cout(\counter_comb_bita4~COUT ),
	.shareout());
defparam counter_comb_bita4.extended_lut = "off";
defparam counter_comb_bita4.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita4.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita5(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita4~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita5~sumout ),
	.cout(),
	.shareout());
defparam counter_comb_bita5.extended_lut = "off";
defparam counter_comb_bita5.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita5.shared_arith = "off";

endmodule

module first_nios2_system_cntr_jgb_1 (
	r_sync_rst,
	wr_rfifo,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	counter_reg_bit_5,
	clock)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
input 	wr_rfifo;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
output 	counter_reg_bit_5;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~sumout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~sumout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~sumout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~sumout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~sumout ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~sumout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wr_rfifo),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wr_rfifo),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wr_rfifo),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wr_rfifo),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wr_rfifo),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wr_rfifo),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

cyclonev_lcell_comb counter_comb_bita0(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita0~sumout ),
	.cout(\counter_comb_bita0~COUT ),
	.shareout());
defparam counter_comb_bita0.extended_lut = "off";
defparam counter_comb_bita0.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita0.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita1(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita0~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita1~sumout ),
	.cout(\counter_comb_bita1~COUT ),
	.shareout());
defparam counter_comb_bita1.extended_lut = "off";
defparam counter_comb_bita1.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita1.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita2(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita1~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita2~sumout ),
	.cout(\counter_comb_bita2~COUT ),
	.shareout());
defparam counter_comb_bita2.extended_lut = "off";
defparam counter_comb_bita2.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita2.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita3(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita2~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita3~sumout ),
	.cout(\counter_comb_bita3~COUT ),
	.shareout());
defparam counter_comb_bita3.extended_lut = "off";
defparam counter_comb_bita3.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita3.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita4(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita3~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita4~sumout ),
	.cout(\counter_comb_bita4~COUT ),
	.shareout());
defparam counter_comb_bita4.extended_lut = "off";
defparam counter_comb_bita4.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita4.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita5(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita4~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita5~sumout ),
	.cout(),
	.shareout());
defparam counter_comb_bita5.extended_lut = "off";
defparam counter_comb_bita5.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita5.shared_arith = "off";

endmodule

module first_nios2_system_first_nios2_system_jtag_uart_scfifo_w (
	q_b_7,
	q_b_0,
	q_b_1,
	q_b_2,
	q_b_3,
	q_b_4,
	q_b_5,
	q_b_6,
	A_st_data_0,
	r_sync_rst,
	A_st_data_1,
	A_st_data_2,
	A_st_data_3,
	A_st_data_4,
	A_st_data_5,
	A_st_data_6,
	A_st_data_7,
	b_full,
	counter_reg_bit_3,
	counter_reg_bit_0,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_5,
	counter_reg_bit_4,
	fifo_wr,
	rvalid0,
	b_non_empty,
	r_val,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_7;
output 	q_b_0;
output 	q_b_1;
output 	q_b_2;
output 	q_b_3;
output 	q_b_4;
output 	q_b_5;
output 	q_b_6;
input 	A_st_data_0;
input 	r_sync_rst;
input 	A_st_data_1;
input 	A_st_data_2;
input 	A_st_data_3;
input 	A_st_data_4;
input 	A_st_data_5;
input 	A_st_data_6;
input 	A_st_data_7;
output 	b_full;
output 	counter_reg_bit_3;
output 	counter_reg_bit_0;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
input 	fifo_wr;
input 	rvalid0;
output 	b_non_empty;
input 	r_val;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



first_nios2_system_scfifo_2 wfifo(
	.q({q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.data({A_st_data_7,A_st_data_6,A_st_data_5,A_st_data_4,A_st_data_3,A_st_data_2,A_st_data_1,A_st_data_0}),
	.r_sync_rst(r_sync_rst),
	.b_full(b_full),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.wrreq(fifo_wr),
	.rvalid0(rvalid0),
	.b_non_empty(b_non_empty),
	.r_val(r_val),
	.clock(clk_clk));

endmodule

module first_nios2_system_scfifo_2 (
	q,
	data,
	r_sync_rst,
	b_full,
	counter_reg_bit_3,
	counter_reg_bit_0,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_5,
	counter_reg_bit_4,
	wrreq,
	rvalid0,
	b_non_empty,
	r_val,
	clock)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q;
input 	[7:0] data;
input 	r_sync_rst;
output 	b_full;
output 	counter_reg_bit_3;
output 	counter_reg_bit_0;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
input 	wrreq;
input 	rvalid0;
output 	b_non_empty;
input 	r_val;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



first_nios2_system_scfifo_3291_1 auto_generated(
	.q({q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.data({data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.r_sync_rst(r_sync_rst),
	.b_full(b_full),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.wrreq(wrreq),
	.rvalid0(rvalid0),
	.b_non_empty(b_non_empty),
	.r_val(r_val),
	.clock(clock));

endmodule

module first_nios2_system_scfifo_3291_1 (
	q,
	data,
	r_sync_rst,
	b_full,
	counter_reg_bit_3,
	counter_reg_bit_0,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_5,
	counter_reg_bit_4,
	wrreq,
	rvalid0,
	b_non_empty,
	r_val,
	clock)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q;
input 	[7:0] data;
input 	r_sync_rst;
output 	b_full;
output 	counter_reg_bit_3;
output 	counter_reg_bit_0;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
input 	wrreq;
input 	rvalid0;
output 	b_non_empty;
input 	r_val;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



first_nios2_system_a_dpfifo_5771_1 dpfifo(
	.q({q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.data({data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.r_sync_rst(r_sync_rst),
	.b_full(b_full),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.wreq(wrreq),
	.rvalid0(rvalid0),
	.b_non_empty(b_non_empty),
	.r_val(r_val),
	.clock(clock));

endmodule

module first_nios2_system_a_dpfifo_5771_1 (
	q,
	data,
	r_sync_rst,
	b_full,
	counter_reg_bit_3,
	counter_reg_bit_0,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_5,
	counter_reg_bit_4,
	wreq,
	rvalid0,
	b_non_empty,
	r_val,
	clock)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q;
input 	[7:0] data;
input 	r_sync_rst;
output 	b_full;
output 	counter_reg_bit_3;
output 	counter_reg_bit_0;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
input 	wreq;
input 	rvalid0;
output 	b_non_empty;
input 	r_val;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wr_ptr|counter_reg_bit[0]~q ;
wire \wr_ptr|counter_reg_bit[1]~q ;
wire \wr_ptr|counter_reg_bit[2]~q ;
wire \wr_ptr|counter_reg_bit[3]~q ;
wire \wr_ptr|counter_reg_bit[4]~q ;
wire \wr_ptr|counter_reg_bit[5]~q ;
wire \rd_ptr_count|counter_reg_bit[0]~q ;
wire \rd_ptr_count|counter_reg_bit[1]~q ;
wire \rd_ptr_count|counter_reg_bit[2]~q ;
wire \rd_ptr_count|counter_reg_bit[3]~q ;
wire \rd_ptr_count|counter_reg_bit[4]~q ;
wire \rd_ptr_count|counter_reg_bit[5]~q ;


first_nios2_system_cntr_jgb_3 wr_ptr(
	.r_sync_rst(r_sync_rst),
	.fifo_wr(wreq),
	.counter_reg_bit_0(\wr_ptr|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\wr_ptr|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\wr_ptr|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\wr_ptr|counter_reg_bit[3]~q ),
	.counter_reg_bit_4(\wr_ptr|counter_reg_bit[4]~q ),
	.counter_reg_bit_5(\wr_ptr|counter_reg_bit[5]~q ),
	.clock(clock));

first_nios2_system_cntr_jgb_2 rd_ptr_count(
	.r_sync_rst(r_sync_rst),
	.r_val(r_val),
	.counter_reg_bit_0(\rd_ptr_count|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\rd_ptr_count|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\rd_ptr_count|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\rd_ptr_count|counter_reg_bit[3]~q ),
	.counter_reg_bit_4(\rd_ptr_count|counter_reg_bit[4]~q ),
	.counter_reg_bit_5(\rd_ptr_count|counter_reg_bit[5]~q ),
	.clock(clock));

first_nios2_system_altsyncram_7pu1_1 FIFOram(
	.q_b({q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.data_a({data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.wren_a(wreq),
	.clocken1(r_val),
	.address_a({\wr_ptr|counter_reg_bit[5]~q ,\wr_ptr|counter_reg_bit[4]~q ,\wr_ptr|counter_reg_bit[3]~q ,\wr_ptr|counter_reg_bit[2]~q ,\wr_ptr|counter_reg_bit[1]~q ,\wr_ptr|counter_reg_bit[0]~q }),
	.address_b({\rd_ptr_count|counter_reg_bit[5]~q ,\rd_ptr_count|counter_reg_bit[4]~q ,\rd_ptr_count|counter_reg_bit[3]~q ,\rd_ptr_count|counter_reg_bit[2]~q ,\rd_ptr_count|counter_reg_bit[1]~q ,\rd_ptr_count|counter_reg_bit[0]~q }),
	.clock1(clock),
	.clock0(clock));

first_nios2_system_a_fefifo_7cf_1 fifo_state(
	.r_sync_rst(r_sync_rst),
	.b_full1(b_full),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.fifo_wr(wreq),
	.rvalid0(rvalid0),
	.b_non_empty1(b_non_empty),
	.r_val(r_val),
	.clock(clock));

endmodule

module first_nios2_system_a_fefifo_7cf_1 (
	r_sync_rst,
	b_full1,
	counter_reg_bit_3,
	counter_reg_bit_0,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_5,
	counter_reg_bit_4,
	fifo_wr,
	rvalid0,
	b_non_empty1,
	r_val,
	clock)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
output 	b_full1;
output 	counter_reg_bit_3;
output 	counter_reg_bit_0;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
input 	fifo_wr;
input 	rvalid0;
output 	b_non_empty1;
input 	r_val;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \_~0_combout ;
wire \b_full~0_combout ;
wire \b_full~1_combout ;
wire \b_non_empty~0_combout ;
wire \b_non_empty~1_combout ;
wire \b_non_empty~2_combout ;


first_nios2_system_cntr_vg7_1 count_usedw(
	.r_sync_rst(r_sync_rst),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.fifo_wr(fifo_wr),
	._(\_~0_combout ),
	.clock(clock));

cyclonev_lcell_comb \_~0 (
	.dataa(!rvalid0),
	.datab(!fifo_wr),
	.datac(!b_non_empty1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\_~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \_~0 .extended_lut = "off";
defparam \_~0 .lut_mask = 64'h9696969696969696;
defparam \_~0 .shared_arith = "off";

dffeas b_full(
	.clk(clock),
	.d(\b_full~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(b_full1),
	.prn(vcc));
defparam b_full.is_wysiwyg = "true";
defparam b_full.power_up = "low";

dffeas b_non_empty(
	.clk(clock),
	.d(\b_non_empty~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(b_non_empty1),
	.prn(vcc));
defparam b_non_empty.is_wysiwyg = "true";
defparam b_non_empty.power_up = "low";

cyclonev_lcell_comb \b_full~0 (
	.dataa(!counter_reg_bit_3),
	.datab(!counter_reg_bit_5),
	.datac(!counter_reg_bit_4),
	.datad(!fifo_wr),
	.datae(!b_non_empty1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\b_full~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \b_full~0 .extended_lut = "off";
defparam \b_full~0 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \b_full~0 .shared_arith = "off";

cyclonev_lcell_comb \b_full~1 (
	.dataa(!b_full1),
	.datab(!counter_reg_bit_0),
	.datac(!counter_reg_bit_2),
	.datad(!counter_reg_bit_1),
	.datae(!r_val),
	.dataf(!\b_full~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\b_full~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \b_full~1 .extended_lut = "off";
defparam \b_full~1 .lut_mask = 64'hFFFF7FFFFFFFFFFF;
defparam \b_full~1 .shared_arith = "off";

cyclonev_lcell_comb \b_non_empty~0 (
	.dataa(!counter_reg_bit_2),
	.datab(!counter_reg_bit_1),
	.datac(!counter_reg_bit_5),
	.datad(!counter_reg_bit_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\b_non_empty~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \b_non_empty~0 .extended_lut = "off";
defparam \b_non_empty~0 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \b_non_empty~0 .shared_arith = "off";

cyclonev_lcell_comb \b_non_empty~1 (
	.dataa(!rvalid0),
	.datab(!counter_reg_bit_3),
	.datac(!counter_reg_bit_0),
	.datad(!b_non_empty1),
	.datae(!\b_non_empty~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\b_non_empty~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \b_non_empty~1 .extended_lut = "off";
defparam \b_non_empty~1 .lut_mask = 64'hFFFFFBFFFFFFFBFF;
defparam \b_non_empty~1 .shared_arith = "off";

cyclonev_lcell_comb \b_non_empty~2 (
	.dataa(!b_full1),
	.datab(!fifo_wr),
	.datac(!\b_non_empty~1_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\b_non_empty~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \b_non_empty~2 .extended_lut = "off";
defparam \b_non_empty~2 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \b_non_empty~2 .shared_arith = "off";

endmodule

module first_nios2_system_cntr_vg7_1 (
	r_sync_rst,
	counter_reg_bit_3,
	counter_reg_bit_0,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_5,
	counter_reg_bit_4,
	fifo_wr,
	_,
	clock)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
output 	counter_reg_bit_3;
output 	counter_reg_bit_0;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
input 	fifo_wr;
input 	_;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~sumout ;
wire \counter_comb_bita0~sumout ;
wire \counter_comb_bita2~sumout ;
wire \counter_comb_bita1~sumout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~sumout ;
wire \counter_comb_bita4~sumout ;


dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

cyclonev_lcell_comb counter_comb_bita0(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita0~sumout ),
	.cout(\counter_comb_bita0~COUT ),
	.shareout());
defparam counter_comb_bita0.extended_lut = "off";
defparam counter_comb_bita0.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita0.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita1(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_1),
	.datae(gnd),
	.dataf(!fifo_wr),
	.datag(gnd),
	.cin(\counter_comb_bita0~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita1~sumout ),
	.cout(\counter_comb_bita1~COUT ),
	.shareout());
defparam counter_comb_bita1.extended_lut = "off";
defparam counter_comb_bita1.lut_mask = 64'h000000FF000000FF;
defparam counter_comb_bita1.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita2(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_2),
	.datae(gnd),
	.dataf(!fifo_wr),
	.datag(gnd),
	.cin(\counter_comb_bita1~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita2~sumout ),
	.cout(\counter_comb_bita2~COUT ),
	.shareout());
defparam counter_comb_bita2.extended_lut = "off";
defparam counter_comb_bita2.lut_mask = 64'h000000FF000000FF;
defparam counter_comb_bita2.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita3(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_3),
	.datae(gnd),
	.dataf(!fifo_wr),
	.datag(gnd),
	.cin(\counter_comb_bita2~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita3~sumout ),
	.cout(\counter_comb_bita3~COUT ),
	.shareout());
defparam counter_comb_bita3.extended_lut = "off";
defparam counter_comb_bita3.lut_mask = 64'h000000FF000000FF;
defparam counter_comb_bita3.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita4(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_4),
	.datae(gnd),
	.dataf(!fifo_wr),
	.datag(gnd),
	.cin(\counter_comb_bita3~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita4~sumout ),
	.cout(\counter_comb_bita4~COUT ),
	.shareout());
defparam counter_comb_bita4.extended_lut = "off";
defparam counter_comb_bita4.lut_mask = 64'h000000FF000000FF;
defparam counter_comb_bita4.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita5(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_5),
	.datae(gnd),
	.dataf(!fifo_wr),
	.datag(gnd),
	.cin(\counter_comb_bita4~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita5~sumout ),
	.cout(),
	.shareout());
defparam counter_comb_bita5.extended_lut = "off";
defparam counter_comb_bita5.lut_mask = 64'h000000FF000000FF;
defparam counter_comb_bita5.shared_arith = "off";

endmodule

module first_nios2_system_altsyncram_7pu1_1 (
	q_b,
	data_a,
	wren_a,
	clocken1,
	address_a,
	address_b,
	clock1,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q_b;
input 	[7:0] data_a;
input 	wren_a;
input 	clocken1;
input 	[5:0] address_a;
input 	[5:0] address_b;
input 	clock1;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

cyclonev_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk1_core_clock_enable = "ena1";
defparam ram_block1a7.clk1_input_clock_enable = "ena1";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "first_nios2_system_jtag_uart:jtag_uart|first_nios2_system_jtag_uart_scfifo_w:the_first_nios2_system_jtag_uart_scfifo_w|scfifo:wfifo|scfifo_3291:auto_generated|a_dpfifo_5771:dpfifo|altsyncram_7pu1:FIFOram|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 6;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 63;
defparam ram_block1a7.port_a_logical_ram_depth = 64;
defparam ram_block1a7.port_a_logical_ram_width = 8;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 6;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "none";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 63;
defparam ram_block1a7.port_b_logical_ram_depth = 64;
defparam ram_block1a7.port_b_logical_ram_width = 8;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";

cyclonev_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk1_core_clock_enable = "ena1";
defparam ram_block1a0.clk1_input_clock_enable = "ena1";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "first_nios2_system_jtag_uart:jtag_uart|first_nios2_system_jtag_uart_scfifo_w:the_first_nios2_system_jtag_uart_scfifo_w|scfifo:wfifo|scfifo_3291:auto_generated|a_dpfifo_5771:dpfifo|altsyncram_7pu1:FIFOram|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 6;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 63;
defparam ram_block1a0.port_a_logical_ram_depth = 64;
defparam ram_block1a0.port_a_logical_ram_width = 8;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock1";
defparam ram_block1a0.port_b_address_width = 6;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "none";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 63;
defparam ram_block1a0.port_b_logical_ram_depth = 64;
defparam ram_block1a0.port_b_logical_ram_width = 8;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock1";
defparam ram_block1a0.ram_block_type = "auto";

cyclonev_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk1_core_clock_enable = "ena1";
defparam ram_block1a1.clk1_input_clock_enable = "ena1";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "first_nios2_system_jtag_uart:jtag_uart|first_nios2_system_jtag_uart_scfifo_w:the_first_nios2_system_jtag_uart_scfifo_w|scfifo:wfifo|scfifo_3291:auto_generated|a_dpfifo_5771:dpfifo|altsyncram_7pu1:FIFOram|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 6;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 63;
defparam ram_block1a1.port_a_logical_ram_depth = 64;
defparam ram_block1a1.port_a_logical_ram_width = 8;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock1";
defparam ram_block1a1.port_b_address_width = 6;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "none";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 63;
defparam ram_block1a1.port_b_logical_ram_depth = 64;
defparam ram_block1a1.port_b_logical_ram_width = 8;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock1";
defparam ram_block1a1.ram_block_type = "auto";

cyclonev_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk1_core_clock_enable = "ena1";
defparam ram_block1a2.clk1_input_clock_enable = "ena1";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "first_nios2_system_jtag_uart:jtag_uart|first_nios2_system_jtag_uart_scfifo_w:the_first_nios2_system_jtag_uart_scfifo_w|scfifo:wfifo|scfifo_3291:auto_generated|a_dpfifo_5771:dpfifo|altsyncram_7pu1:FIFOram|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 6;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 63;
defparam ram_block1a2.port_a_logical_ram_depth = 64;
defparam ram_block1a2.port_a_logical_ram_width = 8;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock1";
defparam ram_block1a2.port_b_address_width = 6;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "none";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 63;
defparam ram_block1a2.port_b_logical_ram_depth = 64;
defparam ram_block1a2.port_b_logical_ram_width = 8;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock1";
defparam ram_block1a2.ram_block_type = "auto";

cyclonev_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk1_core_clock_enable = "ena1";
defparam ram_block1a3.clk1_input_clock_enable = "ena1";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "first_nios2_system_jtag_uart:jtag_uart|first_nios2_system_jtag_uart_scfifo_w:the_first_nios2_system_jtag_uart_scfifo_w|scfifo:wfifo|scfifo_3291:auto_generated|a_dpfifo_5771:dpfifo|altsyncram_7pu1:FIFOram|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 6;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 63;
defparam ram_block1a3.port_a_logical_ram_depth = 64;
defparam ram_block1a3.port_a_logical_ram_width = 8;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock1";
defparam ram_block1a3.port_b_address_width = 6;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "none";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 63;
defparam ram_block1a3.port_b_logical_ram_depth = 64;
defparam ram_block1a3.port_b_logical_ram_width = 8;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock1";
defparam ram_block1a3.ram_block_type = "auto";

cyclonev_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk1_core_clock_enable = "ena1";
defparam ram_block1a4.clk1_input_clock_enable = "ena1";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "first_nios2_system_jtag_uart:jtag_uart|first_nios2_system_jtag_uart_scfifo_w:the_first_nios2_system_jtag_uart_scfifo_w|scfifo:wfifo|scfifo_3291:auto_generated|a_dpfifo_5771:dpfifo|altsyncram_7pu1:FIFOram|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 6;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 63;
defparam ram_block1a4.port_a_logical_ram_depth = 64;
defparam ram_block1a4.port_a_logical_ram_width = 8;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock1";
defparam ram_block1a4.port_b_address_width = 6;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "none";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 63;
defparam ram_block1a4.port_b_logical_ram_depth = 64;
defparam ram_block1a4.port_b_logical_ram_width = 8;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock1";
defparam ram_block1a4.ram_block_type = "auto";

cyclonev_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk1_core_clock_enable = "ena1";
defparam ram_block1a5.clk1_input_clock_enable = "ena1";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "first_nios2_system_jtag_uart:jtag_uart|first_nios2_system_jtag_uart_scfifo_w:the_first_nios2_system_jtag_uart_scfifo_w|scfifo:wfifo|scfifo_3291:auto_generated|a_dpfifo_5771:dpfifo|altsyncram_7pu1:FIFOram|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 6;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 63;
defparam ram_block1a5.port_a_logical_ram_depth = 64;
defparam ram_block1a5.port_a_logical_ram_width = 8;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 6;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "none";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 63;
defparam ram_block1a5.port_b_logical_ram_depth = 64;
defparam ram_block1a5.port_b_logical_ram_width = 8;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";

cyclonev_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk1_core_clock_enable = "ena1";
defparam ram_block1a6.clk1_input_clock_enable = "ena1";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "first_nios2_system_jtag_uart:jtag_uart|first_nios2_system_jtag_uart_scfifo_w:the_first_nios2_system_jtag_uart_scfifo_w|scfifo:wfifo|scfifo_3291:auto_generated|a_dpfifo_5771:dpfifo|altsyncram_7pu1:FIFOram|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 6;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 63;
defparam ram_block1a6.port_a_logical_ram_depth = 64;
defparam ram_block1a6.port_a_logical_ram_width = 8;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 6;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "none";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 63;
defparam ram_block1a6.port_b_logical_ram_depth = 64;
defparam ram_block1a6.port_b_logical_ram_width = 8;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";

endmodule

module first_nios2_system_cntr_jgb_2 (
	r_sync_rst,
	r_val,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	counter_reg_bit_5,
	clock)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
input 	r_val;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
output 	counter_reg_bit_5;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~sumout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~sumout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~sumout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~sumout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~sumout ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~sumout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(r_val),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(r_val),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(r_val),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(r_val),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(r_val),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(r_val),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

cyclonev_lcell_comb counter_comb_bita0(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita0~sumout ),
	.cout(\counter_comb_bita0~COUT ),
	.shareout());
defparam counter_comb_bita0.extended_lut = "off";
defparam counter_comb_bita0.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita0.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita1(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita0~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita1~sumout ),
	.cout(\counter_comb_bita1~COUT ),
	.shareout());
defparam counter_comb_bita1.extended_lut = "off";
defparam counter_comb_bita1.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita1.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita2(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita1~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita2~sumout ),
	.cout(\counter_comb_bita2~COUT ),
	.shareout());
defparam counter_comb_bita2.extended_lut = "off";
defparam counter_comb_bita2.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita2.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita3(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita2~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita3~sumout ),
	.cout(\counter_comb_bita3~COUT ),
	.shareout());
defparam counter_comb_bita3.extended_lut = "off";
defparam counter_comb_bita3.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita3.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita4(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita3~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita4~sumout ),
	.cout(\counter_comb_bita4~COUT ),
	.shareout());
defparam counter_comb_bita4.extended_lut = "off";
defparam counter_comb_bita4.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita4.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita5(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita4~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita5~sumout ),
	.cout(),
	.shareout());
defparam counter_comb_bita5.extended_lut = "off";
defparam counter_comb_bita5.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita5.shared_arith = "off";

endmodule

module first_nios2_system_cntr_jgb_3 (
	r_sync_rst,
	fifo_wr,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	counter_reg_bit_5,
	clock)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
input 	fifo_wr;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
output 	counter_reg_bit_5;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~sumout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~sumout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~sumout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~sumout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~sumout ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~sumout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_wr),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_wr),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_wr),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_wr),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_wr),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_wr),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

cyclonev_lcell_comb counter_comb_bita0(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita0~sumout ),
	.cout(\counter_comb_bita0~COUT ),
	.shareout());
defparam counter_comb_bita0.extended_lut = "off";
defparam counter_comb_bita0.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita0.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita1(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita0~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita1~sumout ),
	.cout(\counter_comb_bita1~COUT ),
	.shareout());
defparam counter_comb_bita1.extended_lut = "off";
defparam counter_comb_bita1.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita1.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita2(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita1~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita2~sumout ),
	.cout(\counter_comb_bita2~COUT ),
	.shareout());
defparam counter_comb_bita2.extended_lut = "off";
defparam counter_comb_bita2.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita2.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita3(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita2~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita3~sumout ),
	.cout(\counter_comb_bita3~COUT ),
	.shareout());
defparam counter_comb_bita3.extended_lut = "off";
defparam counter_comb_bita3.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita3.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita4(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita3~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita4~sumout ),
	.cout(\counter_comb_bita4~COUT ),
	.shareout());
defparam counter_comb_bita4.extended_lut = "off";
defparam counter_comb_bita4.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita4.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita5(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita4~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita5~sumout ),
	.cout(),
	.shareout());
defparam counter_comb_bita5.extended_lut = "off";
defparam counter_comb_bita5.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita5.shared_arith = "off";

endmodule

module first_nios2_system_first_nios2_system_leds (
	data_out_0,
	data_out_1,
	data_out_2,
	data_out_3,
	data_out_4,
	data_out_5,
	data_out_6,
	data_out_7,
	writedata,
	clr_break_line,
	d_write,
	Equal0,
	reset_n,
	wait_latency_counter_1,
	mem_used_1,
	Equal16,
	wait_latency_counter_0,
	clk)/* synthesis synthesis_greybox=1 */;
output 	data_out_0;
output 	data_out_1;
output 	data_out_2;
output 	data_out_3;
output 	data_out_4;
output 	data_out_5;
output 	data_out_6;
output 	data_out_7;
input 	[31:0] writedata;
input 	clr_break_line;
input 	d_write;
input 	Equal0;
input 	reset_n;
input 	wait_latency_counter_1;
input 	mem_used_1;
input 	Equal16;
input 	wait_latency_counter_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \always0~0_combout ;
wire \always0~1_combout ;


dffeas \data_out[0] (
	.clk(clk),
	.d(writedata[0]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_0),
	.prn(vcc));
defparam \data_out[0] .is_wysiwyg = "true";
defparam \data_out[0] .power_up = "low";

dffeas \data_out[1] (
	.clk(clk),
	.d(writedata[1]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_1),
	.prn(vcc));
defparam \data_out[1] .is_wysiwyg = "true";
defparam \data_out[1] .power_up = "low";

dffeas \data_out[2] (
	.clk(clk),
	.d(writedata[2]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_2),
	.prn(vcc));
defparam \data_out[2] .is_wysiwyg = "true";
defparam \data_out[2] .power_up = "low";

dffeas \data_out[3] (
	.clk(clk),
	.d(writedata[3]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_3),
	.prn(vcc));
defparam \data_out[3] .is_wysiwyg = "true";
defparam \data_out[3] .power_up = "low";

dffeas \data_out[4] (
	.clk(clk),
	.d(writedata[4]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_4),
	.prn(vcc));
defparam \data_out[4] .is_wysiwyg = "true";
defparam \data_out[4] .power_up = "low";

dffeas \data_out[5] (
	.clk(clk),
	.d(writedata[5]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_5),
	.prn(vcc));
defparam \data_out[5] .is_wysiwyg = "true";
defparam \data_out[5] .power_up = "low";

dffeas \data_out[6] (
	.clk(clk),
	.d(writedata[6]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_6),
	.prn(vcc));
defparam \data_out[6] .is_wysiwyg = "true";
defparam \data_out[6] .power_up = "low";

dffeas \data_out[7] (
	.clk(clk),
	.d(writedata[7]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_7),
	.prn(vcc));
defparam \data_out[7] .is_wysiwyg = "true";
defparam \data_out[7] .power_up = "low";

cyclonev_lcell_comb \always0~0 (
	.dataa(!d_write),
	.datab(!Equal0),
	.datac(!wait_latency_counter_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'hFDFDFDFDFDFDFDFD;
defparam \always0~0 .shared_arith = "off";

cyclonev_lcell_comb \always0~1 (
	.dataa(!clr_break_line),
	.datab(!wait_latency_counter_1),
	.datac(!mem_used_1),
	.datad(!Equal16),
	.datae(!\always0~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~1 .extended_lut = "off";
defparam \always0~1 .lut_mask = 64'hFDFFFFFFFDFFFFFF;
defparam \always0~1 .shared_arith = "off";

endmodule

module first_nios2_system_first_nios2_system_mm_interconnect_0 (
	q_a_0,
	q_a_1,
	q_a_2,
	q_a_3,
	q_a_4,
	q_a_5,
	q_a_6,
	q_a_7,
	av_readdata_pre_22,
	q_a_22,
	q_a_23,
	q_a_24,
	q_a_25,
	q_a_31,
	q_a_21,
	q_a_11,
	q_a_28,
	q_a_10,
	q_a_27,
	q_a_8,
	q_a_9,
	q_a_26,
	av_readdata_pre_20,
	q_a_20,
	av_readdata_pre_19,
	q_a_19,
	q_a_17,
	q_a_30,
	q_a_18,
	q_a_16,
	q_a_15,
	q_a_12,
	q_a_13,
	q_a_14,
	q_a_29,
	readdata_0,
	readdata_01,
	readdata_02,
	readdata_03,
	readdata_04,
	readdata_05,
	readdata_06,
	q_b_0,
	readdata_07,
	readdata_08,
	readdata_1,
	readdata_11,
	readdata_12,
	readdata_13,
	q_b_1,
	readdata_14,
	readdata_15,
	readdata_16,
	readdata_2,
	readdata_21,
	readdata_22,
	readdata_23,
	q_b_2,
	readdata_24,
	readdata_25,
	readdata_26,
	readdata_3,
	readdata_31,
	readdata_32,
	readdata_33,
	readdata_34,
	q_b_3,
	readdata_35,
	readdata_36,
	q_b_4,
	readdata_4,
	readdata_41,
	readdata_42,
	readdata_43,
	readdata_44,
	readdata_5,
	readdata_51,
	readdata_52,
	q_b_5,
	readdata_53,
	readdata_54,
	readdata_6,
	q_b_6,
	readdata_61,
	readdata_62,
	q_b_7,
	readdata_7,
	Add1,
	readdata_221,
	readdata_231,
	readdata_241,
	readdata_251,
	readdata_311,
	readdata_211,
	Add11,
	readdata_111,
	readdata_28,
	readdata_10,
	readdata_27,
	readdata_8,
	readdata_9,
	readdata_261,
	Add12,
	readdata_20,
	Add13,
	readdata_19,
	readdata_17,
	Add14,
	readdata_30,
	readdata_18,
	Add15,
	readdata_161,
	Add16,
	readdata_151,
	readdata_121,
	readdata_131,
	readdata_141,
	readdata_29,
	data_out,
	data_out1,
	data_out_0,
	data_out_1,
	data_out_2,
	data_out_3,
	data_out_4,
	data_out_5,
	data_out_6,
	data_out_01,
	data_out_11,
	data_out_21,
	data_out_31,
	data_out_41,
	data_out_51,
	data_out_61,
	data_out_02,
	data_out_12,
	data_out_22,
	data_out_32,
	data_out_42,
	data_out_52,
	data_out_62,
	data_out_7,
	data_out2,
	A_st_data_0,
	mem_used_1,
	A_mem_baddr_4,
	A_mem_baddr_5,
	A_mem_baddr_8,
	A_mem_baddr_16,
	A_mem_baddr_15,
	A_mem_baddr_14,
	A_mem_baddr_13,
	Equal1,
	A_mem_baddr_12,
	A_mem_baddr_11,
	A_mem_baddr_10,
	A_mem_baddr_9,
	Equal2,
	A_mem_baddr_7,
	A_mem_baddr_6,
	Equal15,
	always0,
	clr_break_line,
	wait_latency_counter_1,
	wait_latency_counter_0,
	d_write,
	A_mem_baddr_3,
	A_mem_baddr_2,
	Equal0,
	r_sync_rst,
	write,
	wait_latency_counter_01,
	wait_latency_counter_11,
	mem_used_11,
	Equal6,
	wait_latency_counter_02,
	A_st_data_1,
	A_st_data_2,
	A_st_data_3,
	A_st_data_4,
	A_st_data_5,
	A_st_data_6,
	wait_latency_counter_12,
	mem_used_12,
	always1,
	wait_latency_counter_03,
	wait_latency_counter_13,
	mem_used_13,
	Equal16,
	wait_latency_counter_04,
	A_st_data_7,
	wait_latency_counter_14,
	m0_write,
	wait_latency_counter_05,
	d_read,
	read_latency_shift_reg,
	cp_valid,
	W_debug_mode,
	read_latency_shift_reg_0,
	WideOr1,
	WideOr11,
	src0_valid,
	src0_valid1,
	read_latency_shift_reg_01,
	WideOr12,
	WideOr13,
	Equal21,
	wait_latency_counter_06,
	mem_used_14,
	wait_latency_counter_15,
	mem_used_15,
	saved_grant_0,
	always11,
	av_waitrequest,
	mem_used_16,
	av_waitrequest1,
	saved_grant_01,
	waitrequest,
	mem_used_17,
	cpu_data_master_waitrequest,
	i_read,
	ic_fill_tag_5,
	ic_fill_tag_4,
	ic_fill_tag_3,
	ic_fill_tag_2,
	ic_fill_tag_1,
	ic_fill_tag_0,
	WideOr14,
	mem,
	WideOr15,
	ien_AE,
	av_readdata_9,
	ien_AF,
	av_readdata_8,
	src_payload,
	ic_fill_ap_offset_0,
	src_data_38,
	ic_fill_line_0,
	src_data_41,
	ic_fill_ap_offset_2,
	src_data_40,
	ic_fill_ap_offset_1,
	src_data_39,
	ic_fill_line_5,
	src_data_46,
	ic_fill_line_4,
	src_data_45,
	ic_fill_line_3,
	src_data_44,
	ic_fill_line_2,
	src_data_43,
	ic_fill_line_1,
	src_data_42,
	src_payload1,
	save_dest_id,
	WideOr0,
	nonposted_cmd_accepted,
	suppress_change_dest_id,
	b_full,
	src_data_0,
	b_full1,
	b_non_empty,
	read_0,
	counter_reg_bit_0,
	src_payload2,
	src_data_1,
	src_data_2,
	src_data_3,
	src_payload3,
	src_payload4,
	src_payload5,
	src_payload6,
	src_payload7,
	A_mem_byte_en_0,
	src_data_32,
	counter_reg_bit_1,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_5,
	av_readdata_pre_221,
	src_payload8,
	av_readdata_pre_23,
	src_payload9,
	av_readdata_pre_24,
	src_payload10,
	av_readdata_pre_25,
	src_payload11,
	av_readdata_pre_31,
	src_payload12,
	av_readdata_pre_21,
	src_payload13,
	src_payload14,
	av_readdata_pre_11,
	src_payload15,
	src_payload16,
	av_readdata_pre_28,
	src_payload17,
	av_readdata_pre_10,
	src_payload18,
	src_payload19,
	av_readdata_pre_27,
	src_payload20,
	av_readdata_pre_8,
	src_payload21,
	src_payload22,
	av_readdata_pre_9,
	src_payload23,
	src_payload24,
	av_readdata_pre_26,
	src_payload25,
	av_readdata_pre_201,
	src_payload26,
	av_readdata_pre_191,
	src_payload27,
	av_readdata_pre_17,
	src_payload28,
	src_payload29,
	av_readdata_pre_30,
	src_payload30,
	av_readdata_pre_18,
	src_payload31,
	src_payload32,
	av_readdata_pre_16,
	src_payload33,
	src_payload34,
	av_readdata_pre_15,
	src_payload35,
	src_payload36,
	av_readdata_pre_12,
	src_payload37,
	src_payload38,
	av_readdata_pre_13,
	src_payload39,
	src_payload40,
	av_readdata_pre_14,
	src_payload41,
	src_payload42,
	av_readdata_pre_29,
	src_payload43,
	src_payload44,
	src_data_381,
	src_data_391,
	src_data_401,
	src_data_411,
	src_data_421,
	src_data_431,
	src_data_441,
	src_data_451,
	src_data_461,
	src_data_47,
	src_data_48,
	src_data_49,
	src_data_50,
	src_data_321,
	readdata_09,
	src_payload45,
	A_st_data_16,
	src_payload46,
	WideOr16,
	src_payload47,
	readdata_110,
	src_payload48,
	readdata_210,
	src_payload49,
	readdata_37,
	readdata_45,
	src_payload50,
	src_payload51,
	readdata_55,
	src_payload52,
	readdata_63,
	src_payload53,
	readdata_71,
	A_st_data_22,
	src_payload54,
	A_mem_byte_en_2,
	src_data_34,
	A_st_data_23,
	src_payload55,
	A_st_data_24,
	src_payload56,
	A_mem_byte_en_3,
	src_data_35,
	A_st_data_25,
	src_payload57,
	A_st_data_31,
	src_payload58,
	A_st_data_21,
	src_payload59,
	A_st_data_11,
	src_payload60,
	A_mem_byte_en_1,
	src_data_33,
	readdata_112,
	A_st_data_28,
	src_payload61,
	A_st_data_10,
	src_payload62,
	ac,
	readdata_101,
	A_st_data_27,
	src_payload63,
	A_st_data_8,
	src_payload64,
	readdata_81,
	A_st_data_9,
	src_payload65,
	readdata_91,
	A_st_data_26,
	src_payload66,
	A_st_data_20,
	src_payload67,
	A_st_data_19,
	src_payload68,
	A_st_data_17,
	src_payload69,
	A_st_data_30,
	src_payload70,
	A_st_data_18,
	src_payload71,
	src_payload72,
	A_st_data_15,
	src_payload73,
	rvalid,
	readdata_152,
	A_st_data_12,
	src_payload74,
	readdata_122,
	A_st_data_13,
	src_payload75,
	readdata_132,
	A_st_data_14,
	src_payload76,
	woverflow,
	readdata_142,
	A_st_data_29,
	src_payload77,
	src_data_26,
	src_data_25,
	src_data_24,
	src_data_23,
	src_data_22,
	src_data_11,
	src_data_01,
	src_data_21,
	src_data_31,
	src_data_4,
	src_data_5,
	src_data_28,
	src_data_311,
	src_data_27,
	src_data_29,
	src_data_30,
	src_data_111,
	src_data_12,
	src_data_13,
	src_data_14,
	src_data_15,
	src_data_16,
	src_payload78,
	src_data_9,
	src_data_211,
	src_data_6,
	src_data_8,
	src_data_17,
	src_data_18,
	src_data_10,
	src_data_7,
	src_data_20,
	src_data_19,
	src_payload79,
	src_data_341,
	src_payload80,
	src_payload81,
	src_payload82,
	src_payload83,
	src_payload84,
	src_payload85,
	src_payload86,
	src_payload87,
	src_payload88,
	src_data_351,
	src_payload89,
	src_payload90,
	src_payload91,
	src_payload92,
	src_payload93,
	src_payload94,
	src_payload95,
	src_data_331,
	src_payload96,
	src_payload97,
	src_payload98,
	src_payload99,
	src_payload100,
	src_payload101,
	src_payload102,
	src_payload103,
	src_payload104,
	src_payload105,
	GND_port,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	q_a_0;
input 	q_a_1;
input 	q_a_2;
input 	q_a_3;
input 	q_a_4;
input 	q_a_5;
input 	q_a_6;
input 	q_a_7;
output 	av_readdata_pre_22;
input 	q_a_22;
input 	q_a_23;
input 	q_a_24;
input 	q_a_25;
input 	q_a_31;
input 	q_a_21;
input 	q_a_11;
input 	q_a_28;
input 	q_a_10;
input 	q_a_27;
input 	q_a_8;
input 	q_a_9;
input 	q_a_26;
output 	av_readdata_pre_20;
input 	q_a_20;
output 	av_readdata_pre_19;
input 	q_a_19;
input 	q_a_17;
input 	q_a_30;
input 	q_a_18;
input 	q_a_16;
input 	q_a_15;
input 	q_a_12;
input 	q_a_13;
input 	q_a_14;
input 	q_a_29;
input 	readdata_0;
input 	readdata_01;
input 	readdata_02;
input 	readdata_03;
input 	readdata_04;
input 	readdata_05;
input 	readdata_06;
input 	q_b_0;
input 	readdata_07;
input 	readdata_08;
input 	readdata_1;
input 	readdata_11;
input 	readdata_12;
input 	readdata_13;
input 	q_b_1;
input 	readdata_14;
input 	readdata_15;
input 	readdata_16;
input 	readdata_2;
input 	readdata_21;
input 	readdata_22;
input 	readdata_23;
input 	q_b_2;
input 	readdata_24;
input 	readdata_25;
input 	readdata_26;
input 	readdata_3;
input 	readdata_31;
input 	readdata_32;
input 	readdata_33;
input 	readdata_34;
input 	q_b_3;
input 	readdata_35;
input 	readdata_36;
input 	q_b_4;
input 	readdata_4;
input 	readdata_41;
input 	readdata_42;
input 	readdata_43;
input 	readdata_44;
input 	readdata_5;
input 	readdata_51;
input 	readdata_52;
input 	q_b_5;
input 	readdata_53;
input 	readdata_54;
input 	readdata_6;
input 	q_b_6;
input 	readdata_61;
input 	readdata_62;
input 	q_b_7;
input 	readdata_7;
input 	Add1;
input 	readdata_221;
input 	readdata_231;
input 	readdata_241;
input 	readdata_251;
input 	readdata_311;
input 	readdata_211;
input 	Add11;
input 	readdata_111;
input 	readdata_28;
input 	readdata_10;
input 	readdata_27;
input 	readdata_8;
input 	readdata_9;
input 	readdata_261;
input 	Add12;
input 	readdata_20;
input 	Add13;
input 	readdata_19;
input 	readdata_17;
input 	Add14;
input 	readdata_30;
input 	readdata_18;
input 	Add15;
input 	readdata_161;
input 	Add16;
input 	readdata_151;
input 	readdata_121;
input 	readdata_131;
input 	readdata_141;
input 	readdata_29;
input 	data_out;
input 	data_out1;
input 	data_out_0;
input 	data_out_1;
input 	data_out_2;
input 	data_out_3;
input 	data_out_4;
input 	data_out_5;
input 	data_out_6;
input 	data_out_01;
input 	data_out_11;
input 	data_out_21;
input 	data_out_31;
input 	data_out_41;
input 	data_out_51;
input 	data_out_61;
input 	data_out_02;
input 	data_out_12;
input 	data_out_22;
input 	data_out_32;
input 	data_out_42;
input 	data_out_52;
input 	data_out_62;
input 	data_out_7;
input 	data_out2;
input 	A_st_data_0;
output 	mem_used_1;
input 	A_mem_baddr_4;
input 	A_mem_baddr_5;
input 	A_mem_baddr_8;
input 	A_mem_baddr_16;
input 	A_mem_baddr_15;
input 	A_mem_baddr_14;
input 	A_mem_baddr_13;
output 	Equal1;
input 	A_mem_baddr_12;
input 	A_mem_baddr_11;
input 	A_mem_baddr_10;
input 	A_mem_baddr_9;
output 	Equal2;
input 	A_mem_baddr_7;
input 	A_mem_baddr_6;
output 	Equal15;
input 	always0;
input 	clr_break_line;
output 	wait_latency_counter_1;
output 	wait_latency_counter_0;
input 	d_write;
input 	A_mem_baddr_3;
input 	A_mem_baddr_2;
input 	Equal0;
input 	r_sync_rst;
output 	write;
output 	wait_latency_counter_01;
output 	wait_latency_counter_11;
output 	mem_used_11;
output 	Equal6;
output 	wait_latency_counter_02;
input 	A_st_data_1;
input 	A_st_data_2;
input 	A_st_data_3;
input 	A_st_data_4;
input 	A_st_data_5;
input 	A_st_data_6;
output 	wait_latency_counter_12;
output 	mem_used_12;
output 	always1;
output 	wait_latency_counter_03;
output 	wait_latency_counter_13;
output 	mem_used_13;
output 	Equal16;
output 	wait_latency_counter_04;
input 	A_st_data_7;
output 	wait_latency_counter_14;
output 	m0_write;
output 	wait_latency_counter_05;
input 	d_read;
output 	read_latency_shift_reg;
output 	cp_valid;
input 	W_debug_mode;
output 	read_latency_shift_reg_0;
output 	WideOr1;
output 	WideOr11;
output 	src0_valid;
output 	src0_valid1;
output 	read_latency_shift_reg_01;
output 	WideOr12;
output 	WideOr13;
output 	Equal21;
output 	wait_latency_counter_06;
output 	mem_used_14;
output 	wait_latency_counter_15;
output 	mem_used_15;
output 	saved_grant_0;
output 	always11;
input 	av_waitrequest;
output 	mem_used_16;
input 	av_waitrequest1;
output 	saved_grant_01;
input 	waitrequest;
output 	mem_used_17;
output 	cpu_data_master_waitrequest;
input 	i_read;
input 	ic_fill_tag_5;
input 	ic_fill_tag_4;
input 	ic_fill_tag_3;
input 	ic_fill_tag_2;
input 	ic_fill_tag_1;
input 	ic_fill_tag_0;
output 	WideOr14;
output 	mem;
output 	WideOr15;
input 	ien_AE;
input 	av_readdata_9;
input 	ien_AF;
input 	av_readdata_8;
output 	src_payload;
input 	ic_fill_ap_offset_0;
output 	src_data_38;
input 	ic_fill_line_0;
output 	src_data_41;
input 	ic_fill_ap_offset_2;
output 	src_data_40;
input 	ic_fill_ap_offset_1;
output 	src_data_39;
input 	ic_fill_line_5;
output 	src_data_46;
input 	ic_fill_line_4;
output 	src_data_45;
input 	ic_fill_line_3;
output 	src_data_44;
input 	ic_fill_line_2;
output 	src_data_43;
input 	ic_fill_line_1;
output 	src_data_42;
output 	src_payload1;
output 	save_dest_id;
output 	WideOr0;
output 	nonposted_cmd_accepted;
output 	suppress_change_dest_id;
input 	b_full;
output 	src_data_0;
input 	b_full1;
input 	b_non_empty;
input 	read_0;
input 	counter_reg_bit_0;
output 	src_payload2;
output 	src_data_1;
output 	src_data_2;
output 	src_data_3;
output 	src_payload3;
output 	src_payload4;
output 	src_payload5;
output 	src_payload6;
output 	src_payload7;
input 	A_mem_byte_en_0;
output 	src_data_32;
input 	counter_reg_bit_1;
input 	counter_reg_bit_4;
input 	counter_reg_bit_3;
input 	counter_reg_bit_2;
input 	counter_reg_bit_5;
output 	av_readdata_pre_221;
output 	src_payload8;
output 	av_readdata_pre_23;
output 	src_payload9;
output 	av_readdata_pre_24;
output 	src_payload10;
output 	av_readdata_pre_25;
output 	src_payload11;
output 	av_readdata_pre_31;
output 	src_payload12;
output 	av_readdata_pre_21;
output 	src_payload13;
output 	src_payload14;
output 	av_readdata_pre_11;
output 	src_payload15;
output 	src_payload16;
output 	av_readdata_pre_28;
output 	src_payload17;
output 	av_readdata_pre_10;
output 	src_payload18;
output 	src_payload19;
output 	av_readdata_pre_27;
output 	src_payload20;
output 	av_readdata_pre_8;
output 	src_payload21;
output 	src_payload22;
output 	av_readdata_pre_9;
output 	src_payload23;
output 	src_payload24;
output 	av_readdata_pre_26;
output 	src_payload25;
output 	av_readdata_pre_201;
output 	src_payload26;
output 	av_readdata_pre_191;
output 	src_payload27;
output 	av_readdata_pre_17;
output 	src_payload28;
output 	src_payload29;
output 	av_readdata_pre_30;
output 	src_payload30;
output 	av_readdata_pre_18;
output 	src_payload31;
output 	src_payload32;
output 	av_readdata_pre_16;
output 	src_payload33;
output 	src_payload34;
output 	av_readdata_pre_15;
output 	src_payload35;
output 	src_payload36;
output 	av_readdata_pre_12;
output 	src_payload37;
output 	src_payload38;
output 	av_readdata_pre_13;
output 	src_payload39;
output 	src_payload40;
output 	av_readdata_pre_14;
output 	src_payload41;
output 	src_payload42;
output 	av_readdata_pre_29;
output 	src_payload43;
output 	src_payload44;
output 	src_data_381;
output 	src_data_391;
output 	src_data_401;
output 	src_data_411;
output 	src_data_421;
output 	src_data_431;
output 	src_data_441;
output 	src_data_451;
output 	src_data_461;
output 	src_data_47;
output 	src_data_48;
output 	src_data_49;
output 	src_data_50;
output 	src_data_321;
input 	readdata_09;
output 	src_payload45;
input 	A_st_data_16;
output 	src_payload46;
output 	WideOr16;
output 	src_payload47;
input 	readdata_110;
output 	src_payload48;
input 	readdata_210;
output 	src_payload49;
input 	readdata_37;
input 	readdata_45;
output 	src_payload50;
output 	src_payload51;
input 	readdata_55;
output 	src_payload52;
input 	readdata_63;
output 	src_payload53;
input 	readdata_71;
input 	A_st_data_22;
output 	src_payload54;
input 	A_mem_byte_en_2;
output 	src_data_34;
input 	A_st_data_23;
output 	src_payload55;
input 	A_st_data_24;
output 	src_payload56;
input 	A_mem_byte_en_3;
output 	src_data_35;
input 	A_st_data_25;
output 	src_payload57;
input 	A_st_data_31;
output 	src_payload58;
input 	A_st_data_21;
output 	src_payload59;
input 	A_st_data_11;
output 	src_payload60;
input 	A_mem_byte_en_1;
output 	src_data_33;
input 	readdata_112;
input 	A_st_data_28;
output 	src_payload61;
input 	A_st_data_10;
output 	src_payload62;
input 	ac;
input 	readdata_101;
input 	A_st_data_27;
output 	src_payload63;
input 	A_st_data_8;
output 	src_payload64;
input 	readdata_81;
input 	A_st_data_9;
output 	src_payload65;
input 	readdata_91;
input 	A_st_data_26;
output 	src_payload66;
input 	A_st_data_20;
output 	src_payload67;
input 	A_st_data_19;
output 	src_payload68;
input 	A_st_data_17;
output 	src_payload69;
input 	A_st_data_30;
output 	src_payload70;
input 	A_st_data_18;
output 	src_payload71;
output 	src_payload72;
input 	A_st_data_15;
output 	src_payload73;
input 	rvalid;
input 	readdata_152;
input 	A_st_data_12;
output 	src_payload74;
input 	readdata_122;
input 	A_st_data_13;
output 	src_payload75;
input 	readdata_132;
input 	A_st_data_14;
output 	src_payload76;
input 	woverflow;
input 	readdata_142;
input 	A_st_data_29;
output 	src_payload77;
output 	src_data_26;
output 	src_data_25;
output 	src_data_24;
output 	src_data_23;
output 	src_data_22;
output 	src_data_11;
output 	src_data_01;
output 	src_data_21;
output 	src_data_31;
output 	src_data_4;
output 	src_data_5;
output 	src_data_28;
output 	src_data_311;
output 	src_data_27;
output 	src_data_29;
output 	src_data_30;
output 	src_data_111;
output 	src_data_12;
output 	src_data_13;
output 	src_data_14;
output 	src_data_15;
output 	src_data_16;
output 	src_payload78;
output 	src_data_9;
output 	src_data_211;
output 	src_data_6;
output 	src_data_8;
output 	src_data_17;
output 	src_data_18;
output 	src_data_10;
output 	src_data_7;
output 	src_data_20;
output 	src_data_19;
output 	src_payload79;
output 	src_data_341;
output 	src_payload80;
output 	src_payload81;
output 	src_payload82;
output 	src_payload83;
output 	src_payload84;
output 	src_payload85;
output 	src_payload86;
output 	src_payload87;
output 	src_payload88;
output 	src_data_351;
output 	src_payload89;
output 	src_payload90;
output 	src_payload91;
output 	src_payload92;
output 	src_payload93;
output 	src_payload94;
output 	src_payload95;
output 	src_data_331;
output 	src_payload96;
output 	src_payload97;
output 	src_payload98;
output 	src_payload99;
output 	src_payload100;
output 	src_payload101;
output 	src_payload102;
output 	src_payload103;
output 	src_payload104;
output 	src_payload105;
input 	GND_port;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \download1_s1_translator|av_readdata_pre[0]~q ;
wire \download2_s1_translator|av_readdata_pre[0]~q ;
wire \hex1_s1_translator|av_readdata_pre[0]~q ;
wire \hex2_s1_translator|av_readdata_pre[0]~q ;
wire \start_s1_translator|av_readdata_pre[0]~q ;
wire \leds_s1_translator|av_readdata_pre[0]~q ;
wire \jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[0]~q ;
wire \leds_s1_translator|av_readdata_pre[1]~q ;
wire \jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[1]~q ;
wire \hex1_s1_translator|av_readdata_pre[1]~q ;
wire \hex2_s1_translator|av_readdata_pre[1]~q ;
wire \leds_s1_translator|av_readdata_pre[2]~q ;
wire \jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[2]~q ;
wire \hex1_s1_translator|av_readdata_pre[2]~q ;
wire \hex2_s1_translator|av_readdata_pre[2]~q ;
wire \hex2_s1_translator|av_readdata_pre[3]~q ;
wire \leds_s1_translator|av_readdata_pre[3]~q ;
wire \hex1_s1_translator|av_readdata_pre[3]~q ;
wire \jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[3]~q ;
wire \jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[4]~q ;
wire \leds_s1_translator|av_readdata_pre[4]~q ;
wire \hex1_s1_translator|av_readdata_pre[4]~q ;
wire \hex2_s1_translator|av_readdata_pre[4]~q ;
wire \hex2_s1_translator|av_readdata_pre[5]~q ;
wire \leds_s1_translator|av_readdata_pre[5]~q ;
wire \hex1_s1_translator|av_readdata_pre[5]~q ;
wire \jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[5]~q ;
wire \hex2_s1_translator|av_readdata_pre[6]~q ;
wire \jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[6]~q ;
wire \leds_s1_translator|av_readdata_pre[6]~q ;
wire \hex1_s1_translator|av_readdata_pre[6]~q ;
wire \jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[7]~q ;
wire \leds_s1_translator|av_readdata_pre[7]~q ;
wire \jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[21]~q ;
wire \jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[17]~q ;
wire \jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[18]~q ;
wire \jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[16]~q ;
wire \download2_s1_translator|wait_latency_counter[1]~q ;
wire \download2_s1_agent_rsp_fifo|mem_used[1]~q ;
wire \router|Equal14~0_combout ;
wire \download2_s1_agent|m0_write~0_combout ;
wire \router|Equal6~0_combout ;
wire \router|Equal2~1_combout ;
wire \start_s1_agent_rsp_fifo|mem_used[1]~q ;
wire \download1_s1_translator|read_latency_shift_reg[0]~q ;
wire \cpu_data_master_translator|read_accepted~q ;
wire \tenout2_s1_agent|m0_write~0_combout ;
wire \cpu_data_master_translator|uav_read~0_combout ;
wire \camstate2_s1_translator|read_latency_shift_reg[0]~q ;
wire \hex1_s1_translator|read_latency_shift_reg[0]~q ;
wire \hex2_s1_translator|read_latency_shift_reg[0]~q ;
wire \tenout1_s1_translator|read_latency_shift_reg[0]~q ;
wire \tenout2_s1_translator|read_latency_shift_reg[0]~q ;
wire \camdata1_s1_translator|read_latency_shift_reg[0]~q ;
wire \camdata2_s1_translator|read_latency_shift_reg[0]~q ;
wire \rtd1_s1_translator|read_latency_shift_reg[0]~q ;
wire \rtd2_s1_translator|read_latency_shift_reg[0]~q ;
wire \start_s1_translator|read_latency_shift_reg[0]~q ;
wire \download2_s1_translator|read_latency_shift_reg[0]~q ;
wire \cpu_debug_mem_slave_translator|read_latency_shift_reg[0]~q ;
wire \cpu_debug_mem_slave_agent_rsp_fifo|mem[0][74]~q ;
wire \cpu_debug_mem_slave_agent_rsp_fifo|mem[0][56]~q ;
wire \onchip_mem_s1_translator|read_latency_shift_reg[0]~q ;
wire \onchip_mem_s1_agent_rsp_fifo|mem[0][74]~q ;
wire \onchip_mem_s1_agent_rsp_fifo|mem[0][56]~q ;
wire \sysid_control_slave_translator|read_latency_shift_reg[0]~q ;
wire \sys_clk_timer_s1_translator|read_latency_shift_reg[0]~q ;
wire \leds_s1_translator|read_latency_shift_reg[0]~q ;
wire \hex1_s1_agent_rsp_fifo|write~0_combout ;
wire \hex2_s1_agent_rsp_fifo|write~0_combout ;
wire \sys_clk_timer_s1_agent_rsp_fifo|write~0_combout ;
wire \router|always1~1_combout ;
wire \router|src_channel[2]~2_combout ;
wire \router|src_channel[2]~3_combout ;
wire \router|Equal1~1_combout ;
wire \download1_s1_agent_rsp_fifo|write~1_combout ;
wire \leds_s1_agent_rsp_fifo|write~0_combout ;
wire \cmd_demux|WideOr0~3_combout ;
wire \camdata1_s1_agent_rsp_fifo|mem_used[1]~q ;
wire \camdata1_s1_translator|wait_latency_counter[1]~q ;
wire \camdata1_s1_translator|wait_latency_counter[0]~q ;
wire \router|always1~3_combout ;
wire \cmd_demux|sink_ready~0_combout ;
wire \router|always1~4_combout ;
wire \tenout1_s1_agent_rsp_fifo|mem_used[1]~q ;
wire \tenout1_s1_translator|wait_latency_counter[1]~q ;
wire \tenout1_s1_translator|wait_latency_counter[0]~q ;
wire \cmd_demux|sink_ready~1_combout ;
wire \router|always1~5_combout ;
wire \tenout2_s1_agent_rsp_fifo|mem_used[1]~q ;
wire \tenout2_s1_translator|wait_latency_counter[1]~q ;
wire \tenout2_s1_translator|wait_latency_counter[0]~q ;
wire \cmd_demux|sink_ready~2_combout ;
wire \camstate1_s1_agent_rsp_fifo|mem_used[1]~q ;
wire \camstate1_s1_translator|av_waitrequest_generated~0_combout ;
wire \cmd_demux|sink_ready~3_combout ;
wire \camstate2_s1_agent_rsp_fifo|mem_used[1]~q ;
wire \router|always1~6_combout ;
wire \camstate2_s1_translator|av_waitrequest_generated~0_combout ;
wire \cmd_demux|sink_ready~4_combout ;
wire \sysid_control_slave_agent_rsp_fifo|mem_used[1]~q ;
wire \sysid_control_slave_translator|wait_latency_counter[1]~q ;
wire \sysid_control_slave_translator|wait_latency_counter[0]~q ;
wire \router|always1~7_combout ;
wire \cmd_demux|sink_ready~5_combout ;
wire \router|always1~9_combout ;
wire \camdata2_s1_agent_rsp_fifo|mem_used[1]~q ;
wire \camdata2_s1_translator|wait_latency_counter[1]~q ;
wire \camdata2_s1_translator|wait_latency_counter[0]~q ;
wire \cmd_demux|sink_ready~6_combout ;
wire \rtd1_s1_agent_rsp_fifo|mem_used[1]~q ;
wire \rtd1_s1_translator|wait_latency_counter[1]~q ;
wire \rtd1_s1_translator|wait_latency_counter[0]~q ;
wire \router|always1~11_combout ;
wire \cmd_demux|sink_ready~7_combout ;
wire \rtd2_s1_agent_rsp_fifo|mem_used[1]~q ;
wire \rtd2_s1_translator|wait_latency_counter[1]~q ;
wire \rtd2_s1_translator|wait_latency_counter[0]~q ;
wire \router|always1~12_combout ;
wire \cmd_demux|sink_ready~8_combout ;
wire \cpu_debug_mem_slave_agent_rsp_fifo|write~0_combout ;
wire \cmd_demux|WideOr0~6_combout ;
wire \hex1_s1_agent|m0_write~0_combout ;
wire \hex1_s1_translator|av_waitrequest_generated~0_combout ;
wire \hex2_s1_agent|m0_write~0_combout ;
wire \hex2_s1_translator|av_waitrequest_generated~0_combout ;
wire \leds_s1_agent|m0_write~0_combout ;
wire \leds_s1_translator|av_waitrequest_generated~0_combout ;
wire \start_s1_translator|av_waitrequest_generated~0_combout ;
wire \download1_s1_translator|read_latency_shift_reg~1_combout ;
wire \cmd_demux|sink_ready~10_combout ;
wire \cmd_demux|sink_ready~11_combout ;
wire \cmd_mux_002|saved_grant[1]~q ;
wire \cpu_instruction_master_limiter|last_dest_id[2]~q ;
wire \cpu_instruction_master_limiter|has_pending_responses~q ;
wire \router_001|Equal1~0_combout ;
wire \cmd_mux_003|saved_grant[1]~q ;
wire \cpu_instruction_master_limiter|last_dest_id[3]~q ;
wire \onchip_mem_s1_agent_rsp_fifo|mem~0_combout ;
wire \onchip_mem_s1_translator|read_latency_shift_reg~0_combout ;
wire \sys_clk_timer_s1_agent|m0_write~0_combout ;
wire \sys_clk_timer_s1_translator|av_waitrequest_generated~0_combout ;
wire \cmd_demux|src3_valid~0_combout ;
wire \cmd_demux_001|src1_valid~0_combout ;
wire \cmd_demux|sink_ready~12_combout ;
wire \camdata1_s1_agent|m0_write~0_combout ;
wire \cmd_demux|sink_ready~13_combout ;
wire \tenout1_s1_agent|m0_write~0_combout ;
wire \cmd_demux|sink_ready~14_combout ;
wire \tenout2_s1_agent|m0_write~1_combout ;
wire \camstate1_s1_agent|m0_write~0_combout ;
wire \camstate2_s1_agent|m0_write~0_combout ;
wire \router|always1~13_combout ;
wire \cmd_demux|sink_ready~15_combout ;
wire \cmd_demux|sink_ready~16_combout ;
wire \camdata2_s1_agent|m0_write~0_combout ;
wire \cmd_demux|sink_ready~17_combout ;
wire \rtd1_s1_agent|m0_write~0_combout ;
wire \cmd_demux|sink_ready~18_combout ;
wire \rtd2_s1_agent|m0_write~0_combout ;
wire \cmd_demux|src2_valid~0_combout ;
wire \cmd_demux_001|src0_valid~0_combout ;
wire \rsp_demux_002|src1_valid~0_combout ;
wire \rsp_demux_003|src1_valid~0_combout ;
wire \cpu_debug_mem_slave_agent_rsp_fifo|mem[0][61]~q ;
wire \onchip_mem_s1_agent_rsp_fifo|mem[0][61]~q ;
wire \cpu_debug_mem_slave_translator|av_readdata_pre[0]~q ;
wire \camstate2_s1_translator|av_readdata_pre[0]~q ;
wire \tenout1_s1_translator|av_readdata_pre[0]~q ;
wire \tenout2_s1_translator|av_readdata_pre[0]~q ;
wire \camstate1_s1_translator|av_readdata_pre[0]~q ;
wire \rtd2_s1_translator|av_readdata_pre[0]~q ;
wire \rtd1_s1_translator|av_readdata_pre[0]~q ;
wire \sys_clk_timer_s1_translator|av_readdata_pre[0]~q ;
wire \camdata1_s1_translator|av_readdata_pre[0]~q ;
wire \camdata2_s1_translator|av_readdata_pre[0]~q ;
wire \tenout2_s1_translator|av_readdata_pre[1]~q ;
wire \cpu_debug_mem_slave_translator|av_readdata_pre[1]~q ;
wire \camdata1_s1_translator|av_readdata_pre[1]~q ;
wire \camstate2_s1_translator|av_readdata_pre[1]~q ;
wire \sysid_control_slave_translator|av_readdata_pre[30]~q ;
wire \sys_clk_timer_s1_translator|av_readdata_pre[1]~q ;
wire \camdata2_s1_translator|av_readdata_pre[1]~q ;
wire \camstate1_s1_translator|av_readdata_pre[1]~q ;
wire \tenout1_s1_translator|av_readdata_pre[1]~q ;
wire \tenout2_s1_translator|av_readdata_pre[2]~q ;
wire \cpu_debug_mem_slave_translator|av_readdata_pre[2]~q ;
wire \camdata1_s1_translator|av_readdata_pre[2]~q ;
wire \camstate2_s1_translator|av_readdata_pre[2]~q ;
wire \sys_clk_timer_s1_translator|av_readdata_pre[2]~q ;
wire \camdata2_s1_translator|av_readdata_pre[2]~q ;
wire \camstate1_s1_translator|av_readdata_pre[2]~q ;
wire \tenout1_s1_translator|av_readdata_pre[2]~q ;
wire \camdata2_s1_translator|av_readdata_pre[3]~q ;
wire \tenout2_s1_translator|av_readdata_pre[3]~q ;
wire \cpu_debug_mem_slave_translator|av_readdata_pre[3]~q ;
wire \camdata1_s1_translator|av_readdata_pre[3]~q ;
wire \tenout1_s1_translator|av_readdata_pre[3]~q ;
wire \sys_clk_timer_s1_translator|av_readdata_pre[3]~q ;
wire \camstate1_s1_translator|av_readdata_pre[3]~q ;
wire \camstate2_s1_translator|av_readdata_pre[3]~q ;
wire \sys_clk_timer_s1_translator|av_readdata_pre[4]~q ;
wire \cpu_debug_mem_slave_translator|av_readdata_pre[4]~q ;
wire \camdata1_s1_translator|av_readdata_pre[4]~q ;
wire \camdata2_s1_translator|av_readdata_pre[4]~q ;
wire \camstate1_s1_translator|av_readdata_pre[4]~q ;
wire \camstate2_s1_translator|av_readdata_pre[4]~q ;
wire \cpu_debug_mem_slave_translator|av_readdata_pre[5]~q ;
wire \camdata1_s1_translator|av_readdata_pre[5]~q ;
wire \camdata2_s1_translator|av_readdata_pre[5]~q ;
wire \sys_clk_timer_s1_translator|av_readdata_pre[5]~q ;
wire \camstate1_s1_translator|av_readdata_pre[5]~q ;
wire \camstate2_s1_translator|av_readdata_pre[5]~q ;
wire \camdata1_s1_translator|av_readdata_pre[6]~q ;
wire \sys_clk_timer_s1_translator|av_readdata_pre[6]~q ;
wire \cpu_debug_mem_slave_translator|av_readdata_pre[6]~q ;
wire \camdata2_s1_translator|av_readdata_pre[6]~q ;
wire \sys_clk_timer_s1_translator|av_readdata_pre[7]~q ;
wire \cpu_debug_mem_slave_translator|av_readdata_pre[7]~q ;
wire \sys_clk_timer_s1_translator|av_readdata_pre[11]~q ;
wire \jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[10]~q ;
wire \sys_clk_timer_s1_translator|av_readdata_pre[10]~q ;
wire \jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[8]~q ;
wire \sys_clk_timer_s1_translator|av_readdata_pre[8]~q ;
wire \jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[9]~q ;
wire \sys_clk_timer_s1_translator|av_readdata_pre[9]~q ;
wire \jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[15]~q ;
wire \sys_clk_timer_s1_translator|av_readdata_pre[15]~q ;
wire \jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[12]~q ;
wire \sys_clk_timer_s1_translator|av_readdata_pre[12]~q ;
wire \jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[13]~q ;
wire \sys_clk_timer_s1_translator|av_readdata_pre[13]~q ;
wire \jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[14]~q ;
wire \sys_clk_timer_s1_translator|av_readdata_pre[14]~q ;


first_nios2_system_altera_merlin_slave_agent_6 download2_s1_agent(
	.A_mem_baddr_5(A_mem_baddr_5),
	.A_mem_baddr_8(A_mem_baddr_8),
	.Equal1(Equal1),
	.Equal2(Equal2),
	.mem_used_1(\download2_s1_agent_rsp_fifo|mem_used[1]~q ),
	.Equal14(\router|Equal14~0_combout ),
	.m0_write(\download2_s1_agent|m0_write~0_combout ));

first_nios2_system_altera_avalon_sc_fifo_5 download1_s1_agent_rsp_fifo(
	.mem_used_1(mem_used_1),
	.Equal15(Equal15),
	.wait_latency_counter_1(wait_latency_counter_1),
	.wait_latency_counter_0(wait_latency_counter_0),
	.reset(r_sync_rst),
	.read_latency_shift_reg_0(\download1_s1_translator|read_latency_shift_reg[0]~q ),
	.m0_write(\tenout2_s1_agent|m0_write~0_combout ),
	.read_latency_shift_reg(read_latency_shift_reg),
	.write(\download1_s1_agent_rsp_fifo|write~1_combout ),
	.read_latency_shift_reg1(\download1_s1_translator|read_latency_shift_reg~1_combout ),
	.clk(clk_clk));

first_nios2_system_altera_avalon_sc_fifo_10 leds_s1_agent_rsp_fifo(
	.reset(r_sync_rst),
	.wait_latency_counter_1(wait_latency_counter_13),
	.mem_used_1(mem_used_13),
	.Equal16(Equal16),
	.wait_latency_counter_0(wait_latency_counter_04),
	.m0_write(\tenout2_s1_agent|m0_write~0_combout ),
	.read_latency_shift_reg(read_latency_shift_reg),
	.read_latency_shift_reg_0(\leds_s1_translator|read_latency_shift_reg[0]~q ),
	.write(\leds_s1_agent_rsp_fifo|write~0_combout ),
	.av_waitrequest_generated(\leds_s1_translator|av_waitrequest_generated~0_combout ),
	.clk(clk_clk));

first_nios2_system_altera_merlin_slave_agent_10 leds_s1_agent(
	.mem_used_1(mem_used_13),
	.Equal16(Equal16),
	.m0_write(\leds_s1_agent|m0_write~0_combout ));

first_nios2_system_altera_avalon_sc_fifo_15 sys_clk_timer_s1_agent_rsp_fifo(
	.reset(r_sync_rst),
	.m0_write(\tenout2_s1_agent|m0_write~0_combout ),
	.read_latency_shift_reg(read_latency_shift_reg),
	.read_latency_shift_reg_0(\sys_clk_timer_s1_translator|read_latency_shift_reg[0]~q ),
	.Equal2(Equal21),
	.wait_latency_counter_0(wait_latency_counter_06),
	.mem_used_1(mem_used_14),
	.wait_latency_counter_1(wait_latency_counter_15),
	.write(\sys_clk_timer_s1_agent_rsp_fifo|write~0_combout ),
	.av_waitrequest_generated(\sys_clk_timer_s1_translator|av_waitrequest_generated~0_combout ),
	.clk(clk_clk));

first_nios2_system_altera_merlin_slave_agent_15 sys_clk_timer_s1_agent(
	.Equal2(Equal21),
	.mem_used_1(mem_used_14),
	.m0_write(\sys_clk_timer_s1_agent|m0_write~0_combout ));

first_nios2_system_altera_avalon_sc_fifo_11 onchip_mem_s1_agent_rsp_fifo(
	.clr_break_line(clr_break_line),
	.reset(r_sync_rst),
	.uav_read(\cpu_data_master_translator|uav_read~0_combout ),
	.read_latency_shift_reg_0(\onchip_mem_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_74_0(\onchip_mem_s1_agent_rsp_fifo|mem[0][74]~q ),
	.mem_56_0(\onchip_mem_s1_agent_rsp_fifo|mem[0][56]~q ),
	.mem_used_1(mem_used_15),
	.saved_grant_0(saved_grant_0),
	.i_read(i_read),
	.saved_grant_1(\cmd_mux_003|saved_grant[1]~q ),
	.WideOr1(WideOr15),
	.mem(\onchip_mem_s1_agent_rsp_fifo|mem~0_combout ),
	.mem_61_0(\onchip_mem_s1_agent_rsp_fifo|mem[0][61]~q ),
	.clk(clk_clk));

first_nios2_system_altera_avalon_sc_fifo_4 cpu_debug_mem_slave_agent_rsp_fifo(
	.reset(r_sync_rst),
	.uav_read(\cpu_data_master_translator|uav_read~0_combout ),
	.read_latency_shift_reg_0(\cpu_debug_mem_slave_translator|read_latency_shift_reg[0]~q ),
	.mem_74_0(\cpu_debug_mem_slave_agent_rsp_fifo|mem[0][74]~q ),
	.mem_56_0(\cpu_debug_mem_slave_agent_rsp_fifo|mem[0][56]~q ),
	.saved_grant_0(saved_grant_01),
	.waitrequest(waitrequest),
	.mem_used_1(mem_used_17),
	.write(\cpu_debug_mem_slave_agent_rsp_fifo|write~0_combout ),
	.saved_grant_1(\cmd_mux_002|saved_grant[1]~q ),
	.i_read(i_read),
	.WideOr1(WideOr14),
	.mem(mem),
	.mem_61_0(\cpu_debug_mem_slave_agent_rsp_fifo|mem[0][61]~q ),
	.clk(clk_clk));

first_nios2_system_altera_avalon_sc_fifo_16 sysid_control_slave_agent_rsp_fifo(
	.reset(r_sync_rst),
	.read_latency_shift_reg_0(\sysid_control_slave_translator|read_latency_shift_reg[0]~q ),
	.mem_used_1(\sysid_control_slave_agent_rsp_fifo|mem_used[1]~q ),
	.sink_ready(\cmd_demux|sink_ready~5_combout ),
	.sink_ready1(\cmd_demux|sink_ready~15_combout ),
	.clk(clk_clk));

first_nios2_system_altera_avalon_sc_fifo_9 jtag_uart_avalon_jtag_slave_agent_rsp_fifo(
	.A_mem_baddr_4(A_mem_baddr_4),
	.A_mem_baddr_3(A_mem_baddr_3),
	.reset(r_sync_rst),
	.read_latency_shift_reg(read_latency_shift_reg),
	.read_latency_shift_reg_0(read_latency_shift_reg_01),
	.av_waitrequest(av_waitrequest),
	.mem_used_1(mem_used_16),
	.always1(\router|always1~13_combout ),
	.clk(clk_clk));

first_nios2_system_altera_merlin_master_agent cpu_data_master_agent(
	.clr_break_line(clr_break_line),
	.d_write(d_write),
	.d_read(d_read),
	.read_accepted(\cpu_data_master_translator|read_accepted~q ),
	.cp_valid(cp_valid));

first_nios2_system_altera_merlin_slave_translator_18 tenout2_s1_translator(
	.av_readdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,readdata_31,readdata_2,readdata_1,readdata_03}),
	.d_write(d_write),
	.reset(r_sync_rst),
	.cp_valid(cp_valid),
	.read_latency_shift_reg_0(\tenout2_s1_translator|read_latency_shift_reg[0]~q ),
	.wait_latency_counter_1(\tenout2_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\tenout2_s1_translator|wait_latency_counter[0]~q ),
	.sink_ready(\cmd_demux|sink_ready~2_combout ),
	.m0_write(\tenout2_s1_agent|m0_write~1_combout ),
	.av_readdata_pre_0(\tenout2_s1_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_1(\tenout2_s1_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_2(\tenout2_s1_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_3(\tenout2_s1_translator|av_readdata_pre[3]~q ),
	.clk(clk_clk));

first_nios2_system_altera_merlin_slave_translator_17 tenout1_s1_translator(
	.av_readdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,readdata_34,readdata_26,readdata_16,readdata_02}),
	.d_write(d_write),
	.reset(r_sync_rst),
	.cp_valid(cp_valid),
	.read_latency_shift_reg_0(\tenout1_s1_translator|read_latency_shift_reg[0]~q ),
	.wait_latency_counter_1(\tenout1_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\tenout1_s1_translator|wait_latency_counter[0]~q ),
	.sink_ready(\cmd_demux|sink_ready~1_combout ),
	.m0_write(\tenout1_s1_agent|m0_write~0_combout ),
	.av_readdata_pre_0(\tenout1_s1_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_1(\tenout1_s1_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_2(\tenout1_s1_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_3(\tenout1_s1_translator|av_readdata_pre[3]~q ),
	.clk(clk_clk));

first_nios2_system_altera_merlin_slave_translator_8 hex2_s1_translator(
	.av_readdata_pre_0(\hex2_s1_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_1(\hex2_s1_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_2(\hex2_s1_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_3(\hex2_s1_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_4(\hex2_s1_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_5(\hex2_s1_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_6(\hex2_s1_translator|av_readdata_pre[6]~q ),
	.av_readdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_out_61,data_out_51,data_out_41,data_out_31,data_out_21,data_out_11,data_out_01}),
	.A_mem_baddr_7(A_mem_baddr_7),
	.clr_break_line(clr_break_line),
	.d_write(d_write),
	.Equal0(Equal0),
	.reset(r_sync_rst),
	.wait_latency_counter_1(wait_latency_counter_12),
	.mem_used_1(mem_used_12),
	.always1(always1),
	.wait_latency_counter_0(wait_latency_counter_03),
	.m0_write(\tenout2_s1_agent|m0_write~0_combout ),
	.uav_read(\cpu_data_master_translator|uav_read~0_combout ),
	.cp_valid(cp_valid),
	.read_latency_shift_reg_0(\hex2_s1_translator|read_latency_shift_reg[0]~q ),
	.m0_write1(\hex2_s1_agent|m0_write~0_combout ),
	.av_waitrequest_generated(\hex2_s1_translator|av_waitrequest_generated~0_combout ),
	.clk(clk_clk));

first_nios2_system_altera_merlin_slave_translator_7 hex1_s1_translator(
	.av_readdata_pre_0(\hex1_s1_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_1(\hex1_s1_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_2(\hex1_s1_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_3(\hex1_s1_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_4(\hex1_s1_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_5(\hex1_s1_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_6(\hex1_s1_translator|av_readdata_pre[6]~q ),
	.av_readdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_out_6,data_out_5,data_out_4,data_out_3,data_out_2,data_out_1,data_out_0}),
	.clr_break_line(clr_break_line),
	.d_write(d_write),
	.Equal0(Equal0),
	.reset(r_sync_rst),
	.wait_latency_counter_1(wait_latency_counter_11),
	.wait_latency_counter_0(wait_latency_counter_02),
	.m0_write(\tenout2_s1_agent|m0_write~0_combout ),
	.uav_read(\cpu_data_master_translator|uav_read~0_combout ),
	.cp_valid(cp_valid),
	.read_latency_shift_reg_0(\hex1_s1_translator|read_latency_shift_reg[0]~q ),
	.m0_write1(\hex1_s1_agent|m0_write~0_combout ),
	.av_waitrequest_generated(\hex1_s1_translator|av_waitrequest_generated~0_combout ),
	.clk(clk_clk));

first_nios2_system_altera_merlin_slave_translator_3 camstate2_s1_translator(
	.av_readdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,readdata_54,readdata_44,readdata_36,readdata_23,readdata_13,readdata_01}),
	.d_write(d_write),
	.reset(r_sync_rst),
	.m0_write(\tenout2_s1_agent|m0_write~0_combout ),
	.cp_valid(cp_valid),
	.read_latency_shift_reg_0(\camstate2_s1_translator|read_latency_shift_reg[0]~q ),
	.always1(\router|always1~1_combout ),
	.mem_used_1(\camstate2_s1_agent_rsp_fifo|mem_used[1]~q ),
	.always11(\router|always1~6_combout ),
	.av_waitrequest_generated(\camstate2_s1_translator|av_waitrequest_generated~0_combout ),
	.sink_ready(\cmd_demux|sink_ready~11_combout ),
	.m0_write1(\camstate2_s1_agent|m0_write~0_combout ),
	.av_readdata_pre_0(\camstate2_s1_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_1(\camstate2_s1_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_2(\camstate2_s1_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_3(\camstate2_s1_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_4(\camstate2_s1_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_5(\camstate2_s1_translator|av_readdata_pre[5]~q ),
	.clk(clk_clk));

first_nios2_system_altera_merlin_slave_translator_2 camstate1_s1_translator(
	.av_readdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,readdata_53,readdata_43,readdata_35,readdata_25,readdata_15,readdata_04}),
	.d_write(d_write),
	.reset(r_sync_rst),
	.Equal6(\router|Equal6~0_combout ),
	.m0_write(\tenout2_s1_agent|m0_write~0_combout ),
	.cp_valid(cp_valid),
	.read_latency_shift_reg_0(read_latency_shift_reg_0),
	.always1(\router|always1~1_combout ),
	.mem_used_1(\camstate1_s1_agent_rsp_fifo|mem_used[1]~q ),
	.av_waitrequest_generated(\camstate1_s1_translator|av_waitrequest_generated~0_combout ),
	.sink_ready(\cmd_demux|sink_ready~10_combout ),
	.m0_write1(\camstate1_s1_agent|m0_write~0_combout ),
	.av_readdata_pre_0(\camstate1_s1_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_1(\camstate1_s1_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_2(\camstate1_s1_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_3(\camstate1_s1_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_4(\camstate1_s1_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_5(\camstate1_s1_translator|av_readdata_pre[5]~q ),
	.clk(clk_clk));

first_nios2_system_altera_merlin_slave_translator_14 start_s1_translator(
	.av_readdata_pre_0(\start_s1_translator|av_readdata_pre[0]~q ),
	.av_readdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_out2}),
	.clr_break_line(clr_break_line),
	.d_write(d_write),
	.Equal0(Equal0),
	.reset(r_sync_rst),
	.wait_latency_counter_1(wait_latency_counter_14),
	.m0_write(m0_write),
	.wait_latency_counter_0(wait_latency_counter_05),
	.m0_write1(\tenout2_s1_agent|m0_write~0_combout ),
	.uav_read(\cpu_data_master_translator|uav_read~0_combout ),
	.cp_valid(cp_valid),
	.read_latency_shift_reg_0(\start_s1_translator|read_latency_shift_reg[0]~q ),
	.av_waitrequest_generated(\start_s1_translator|av_waitrequest_generated~0_combout ),
	.clk(clk_clk));

first_nios2_system_altera_merlin_slave_translator_13 rtd2_s1_translator(
	.av_readdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,readdata_05}),
	.d_write(d_write),
	.reset(r_sync_rst),
	.cp_valid(cp_valid),
	.read_latency_shift_reg_0(\rtd2_s1_translator|read_latency_shift_reg[0]~q ),
	.wait_latency_counter_1(\rtd2_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\rtd2_s1_translator|wait_latency_counter[0]~q ),
	.sink_ready(\cmd_demux|sink_ready~8_combout ),
	.m0_write(\rtd2_s1_agent|m0_write~0_combout ),
	.av_readdata_pre_0(\rtd2_s1_translator|av_readdata_pre[0]~q ),
	.clk(clk_clk));

first_nios2_system_altera_merlin_slave_translator_12 rtd1_s1_translator(
	.av_readdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,readdata_06}),
	.d_write(d_write),
	.reset(r_sync_rst),
	.cp_valid(cp_valid),
	.read_latency_shift_reg_0(\rtd1_s1_translator|read_latency_shift_reg[0]~q ),
	.wait_latency_counter_1(\rtd1_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\rtd1_s1_translator|wait_latency_counter[0]~q ),
	.sink_ready(\cmd_demux|sink_ready~7_combout ),
	.m0_write(\rtd1_s1_agent|m0_write~0_combout ),
	.av_readdata_pre_0(\rtd1_s1_translator|av_readdata_pre[0]~q ),
	.clk(clk_clk));

first_nios2_system_altera_merlin_slave_translator_1 camdata2_s1_translator(
	.av_readdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,readdata_62,readdata_52,readdata_42,readdata_3,readdata_24,readdata_14,readdata_08}),
	.d_write(d_write),
	.reset(r_sync_rst),
	.cp_valid(cp_valid),
	.read_latency_shift_reg_0(\camdata2_s1_translator|read_latency_shift_reg[0]~q ),
	.wait_latency_counter_1(\camdata2_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\camdata2_s1_translator|wait_latency_counter[0]~q ),
	.sink_ready(\cmd_demux|sink_ready~6_combout ),
	.m0_write(\camdata2_s1_agent|m0_write~0_combout ),
	.av_readdata_pre_0(\camdata2_s1_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_1(\camdata2_s1_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_2(\camdata2_s1_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_3(\camdata2_s1_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_4(\camdata2_s1_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_5(\camdata2_s1_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_6(\camdata2_s1_translator|av_readdata_pre[6]~q ),
	.clk(clk_clk));

first_nios2_system_altera_merlin_slave_translator camdata1_s1_translator(
	.av_readdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,readdata_6,readdata_51,readdata_41,readdata_33,readdata_22,readdata_12,readdata_07}),
	.d_write(d_write),
	.reset(r_sync_rst),
	.cp_valid(cp_valid),
	.read_latency_shift_reg_0(\camdata1_s1_translator|read_latency_shift_reg[0]~q ),
	.wait_latency_counter_1(\camdata1_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\camdata1_s1_translator|wait_latency_counter[0]~q ),
	.sink_ready(\cmd_demux|sink_ready~0_combout ),
	.m0_write(\camdata1_s1_agent|m0_write~0_combout ),
	.av_readdata_pre_0(\camdata1_s1_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_1(\camdata1_s1_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_2(\camdata1_s1_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_3(\camdata1_s1_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_4(\camdata1_s1_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_5(\camdata1_s1_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_6(\camdata1_s1_translator|av_readdata_pre[6]~q ),
	.clk(clk_clk));

first_nios2_system_altera_merlin_slave_translator_6 download2_s1_translator(
	.av_readdata_pre_0(\download2_s1_translator|av_readdata_pre[0]~q ),
	.av_readdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_out1}),
	.clr_break_line(clr_break_line),
	.d_write(d_write),
	.Equal0(Equal0),
	.reset(r_sync_rst),
	.wait_latency_counter_1(\download2_s1_translator|wait_latency_counter[1]~q ),
	.m0_write(\download2_s1_agent|m0_write~0_combout ),
	.wait_latency_counter_0(wait_latency_counter_01),
	.uav_read(\cpu_data_master_translator|uav_read~0_combout ),
	.cp_valid(cp_valid),
	.read_latency_shift_reg_0(\download2_s1_translator|read_latency_shift_reg[0]~q ),
	.clk(clk_clk));

first_nios2_system_altera_merlin_slave_translator_5 download1_s1_translator(
	.av_readdata_pre_0(\download1_s1_translator|av_readdata_pre[0]~q ),
	.av_readdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_out}),
	.always0(always0),
	.clr_break_line(clr_break_line),
	.wait_latency_counter_1(wait_latency_counter_1),
	.wait_latency_counter_0(wait_latency_counter_0),
	.d_write(d_write),
	.Equal0(Equal0),
	.reset(r_sync_rst),
	.read_latency_shift_reg_0(\download1_s1_translator|read_latency_shift_reg[0]~q ),
	.uav_read(\cpu_data_master_translator|uav_read~0_combout ),
	.read_latency_shift_reg(read_latency_shift_reg),
	.cp_valid(cp_valid),
	.write(\download1_s1_agent_rsp_fifo|write~1_combout ),
	.read_latency_shift_reg1(\download1_s1_translator|read_latency_shift_reg~1_combout ),
	.clk(clk_clk));

first_nios2_system_altera_merlin_slave_translator_10 leds_s1_translator(
	.av_readdata_pre_0(\leds_s1_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_1(\leds_s1_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_2(\leds_s1_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_3(\leds_s1_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_4(\leds_s1_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_5(\leds_s1_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_6(\leds_s1_translator|av_readdata_pre[6]~q ),
	.av_readdata_pre_7(\leds_s1_translator|av_readdata_pre[7]~q ),
	.av_readdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_out_7,data_out_62,data_out_52,data_out_42,data_out_32,data_out_22,data_out_12,data_out_02}),
	.clr_break_line(clr_break_line),
	.d_write(d_write),
	.Equal0(Equal0),
	.reset(r_sync_rst),
	.wait_latency_counter_1(wait_latency_counter_13),
	.wait_latency_counter_0(wait_latency_counter_04),
	.m0_write(\tenout2_s1_agent|m0_write~0_combout ),
	.uav_read(\cpu_data_master_translator|uav_read~0_combout ),
	.cp_valid(cp_valid),
	.read_latency_shift_reg_0(\leds_s1_translator|read_latency_shift_reg[0]~q ),
	.m0_write1(\leds_s1_agent|m0_write~0_combout ),
	.av_waitrequest_generated(\leds_s1_translator|av_waitrequest_generated~0_combout ),
	.clk(clk_clk));

first_nios2_system_altera_merlin_slave_translator_15 sys_clk_timer_s1_translator(
	.clr_break_line(clr_break_line),
	.d_write(d_write),
	.reset(r_sync_rst),
	.m0_write(\tenout2_s1_agent|m0_write~0_combout ),
	.uav_read(\cpu_data_master_translator|uav_read~0_combout ),
	.cp_valid(cp_valid),
	.read_latency_shift_reg_0(\sys_clk_timer_s1_translator|read_latency_shift_reg[0]~q ),
	.wait_latency_counter_0(wait_latency_counter_06),
	.wait_latency_counter_1(wait_latency_counter_15),
	.m0_write1(\sys_clk_timer_s1_agent|m0_write~0_combout ),
	.av_waitrequest_generated(\sys_clk_timer_s1_translator|av_waitrequest_generated~0_combout ),
	.av_readdata_pre_0(\sys_clk_timer_s1_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_1(\sys_clk_timer_s1_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_2(\sys_clk_timer_s1_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_3(\sys_clk_timer_s1_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_4(\sys_clk_timer_s1_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_5(\sys_clk_timer_s1_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_6(\sys_clk_timer_s1_translator|av_readdata_pre[6]~q ),
	.av_readdata_pre_7(\sys_clk_timer_s1_translator|av_readdata_pre[7]~q ),
	.av_readdata_pre_11(\sys_clk_timer_s1_translator|av_readdata_pre[11]~q ),
	.av_readdata_pre_10(\sys_clk_timer_s1_translator|av_readdata_pre[10]~q ),
	.av_readdata_pre_8(\sys_clk_timer_s1_translator|av_readdata_pre[8]~q ),
	.av_readdata_pre_9(\sys_clk_timer_s1_translator|av_readdata_pre[9]~q ),
	.av_readdata_pre_15(\sys_clk_timer_s1_translator|av_readdata_pre[15]~q ),
	.av_readdata_pre_12(\sys_clk_timer_s1_translator|av_readdata_pre[12]~q ),
	.av_readdata_pre_13(\sys_clk_timer_s1_translator|av_readdata_pre[13]~q ),
	.av_readdata_pre_14(\sys_clk_timer_s1_translator|av_readdata_pre[14]~q ),
	.av_readdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,readdata_152,readdata_142,readdata_132,readdata_122,readdata_112,readdata_101,readdata_91,readdata_81,readdata_71,readdata_63,readdata_55,readdata_45,readdata_37,readdata_210,readdata_110,readdata_09}),
	.clk(clk_clk));

first_nios2_system_altera_merlin_slave_translator_11 onchip_mem_s1_translator(
	.clr_break_line(clr_break_line),
	.reset(r_sync_rst),
	.read_latency_shift_reg_0(\onchip_mem_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_used_1(mem_used_15),
	.WideOr1(WideOr15),
	.mem(\onchip_mem_s1_agent_rsp_fifo|mem~0_combout ),
	.read_latency_shift_reg(\onchip_mem_s1_translator|read_latency_shift_reg~0_combout ),
	.clk(clk_clk));

first_nios2_system_altera_merlin_slave_translator_4 cpu_debug_mem_slave_translator(
	.av_readdata({readdata_311,readdata_30,readdata_29,readdata_28,readdata_27,readdata_261,readdata_251,readdata_241,readdata_231,readdata_221,readdata_211,readdata_20,readdata_19,readdata_18,readdata_17,readdata_161,readdata_151,readdata_141,readdata_131,readdata_121,readdata_111,readdata_10,
readdata_9,readdata_8,readdata_7,readdata_61,readdata_5,readdata_4,readdata_32,readdata_21,readdata_11,readdata_0}),
	.clr_break_line(clr_break_line),
	.reset(r_sync_rst),
	.read_latency_shift_reg_0(\cpu_debug_mem_slave_translator|read_latency_shift_reg[0]~q ),
	.write(\cpu_debug_mem_slave_agent_rsp_fifo|write~0_combout ),
	.WideOr1(WideOr14),
	.mem(mem),
	.av_readdata_pre_0(\cpu_debug_mem_slave_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_1(\cpu_debug_mem_slave_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_2(\cpu_debug_mem_slave_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_3(\cpu_debug_mem_slave_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_4(\cpu_debug_mem_slave_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_5(\cpu_debug_mem_slave_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_6(\cpu_debug_mem_slave_translator|av_readdata_pre[6]~q ),
	.av_readdata_pre_7(\cpu_debug_mem_slave_translator|av_readdata_pre[7]~q ),
	.av_readdata_pre_22(av_readdata_pre_221),
	.av_readdata_pre_23(av_readdata_pre_23),
	.av_readdata_pre_24(av_readdata_pre_24),
	.av_readdata_pre_25(av_readdata_pre_25),
	.av_readdata_pre_31(av_readdata_pre_31),
	.av_readdata_pre_21(av_readdata_pre_21),
	.av_readdata_pre_11(av_readdata_pre_11),
	.av_readdata_pre_28(av_readdata_pre_28),
	.av_readdata_pre_10(av_readdata_pre_10),
	.av_readdata_pre_27(av_readdata_pre_27),
	.av_readdata_pre_8(av_readdata_pre_8),
	.av_readdata_pre_9(av_readdata_pre_9),
	.av_readdata_pre_26(av_readdata_pre_26),
	.av_readdata_pre_20(av_readdata_pre_201),
	.av_readdata_pre_19(av_readdata_pre_191),
	.av_readdata_pre_17(av_readdata_pre_17),
	.av_readdata_pre_30(av_readdata_pre_30),
	.av_readdata_pre_18(av_readdata_pre_18),
	.av_readdata_pre_16(av_readdata_pre_16),
	.av_readdata_pre_15(av_readdata_pre_15),
	.av_readdata_pre_12(av_readdata_pre_12),
	.av_readdata_pre_13(av_readdata_pre_13),
	.av_readdata_pre_14(av_readdata_pre_14),
	.av_readdata_pre_29(av_readdata_pre_29),
	.clk(clk_clk));

first_nios2_system_altera_merlin_slave_translator_16 sysid_control_slave_translator(
	.d_write(d_write),
	.av_readdata({gnd,A_mem_baddr_2,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.reset(r_sync_rst),
	.cp_valid(cp_valid),
	.read_latency_shift_reg_0(\sysid_control_slave_translator|read_latency_shift_reg[0]~q ),
	.mem_used_1(\sysid_control_slave_agent_rsp_fifo|mem_used[1]~q ),
	.wait_latency_counter_1(\sysid_control_slave_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\sysid_control_slave_translator|wait_latency_counter[0]~q ),
	.always1(\router|always1~7_combout ),
	.sink_ready(\cmd_demux|sink_ready~5_combout ),
	.av_readdata_pre_30(\sysid_control_slave_translator|av_readdata_pre[30]~q ),
	.clk(clk_clk));

first_nios2_system_altera_merlin_slave_translator_9 jtag_uart_avalon_jtag_slave_translator(
	.av_readdata_pre_0(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_1(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_2(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_3(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_4(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_5(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_6(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[6]~q ),
	.av_readdata_pre_7(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[7]~q ),
	.av_readdata_pre_22(av_readdata_pre_22),
	.av_readdata_pre_21(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[21]~q ),
	.av_readdata_pre_20(av_readdata_pre_20),
	.av_readdata_pre_19(av_readdata_pre_19),
	.av_readdata_pre_17(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[17]~q ),
	.av_readdata_pre_18(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[18]~q ),
	.av_readdata_pre_16(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[16]~q ),
	.q_b_0(q_b_0),
	.q_b_1(q_b_1),
	.q_b_2(q_b_2),
	.q_b_3(q_b_3),
	.q_b_4(q_b_4),
	.q_b_5(q_b_5),
	.q_b_6(q_b_6),
	.q_b_7(q_b_7),
	.av_readdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,Add1,Add11,Add12,Add13,Add15,Add14,Add16,rvalid,woverflow,gnd,b_non_empty,gnd,ac,av_readdata_9,av_readdata_8,GND_port,GND_port,GND_port,GND_port,GND_port,GND_port,ien_AE,ien_AF}),
	.reset(r_sync_rst),
	.read_latency_shift_reg(read_latency_shift_reg),
	.read_latency_shift_reg_0(read_latency_shift_reg_01),
	.av_waitrequest(av_waitrequest),
	.av_waitrequest1(av_waitrequest1),
	.b_full(b_full),
	.b_full1(b_full1),
	.read_0(read_0),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_5(counter_reg_bit_5),
	.av_readdata_pre_10(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[10]~q ),
	.av_readdata_pre_8(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[8]~q ),
	.av_readdata_pre_9(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[9]~q ),
	.av_readdata_pre_15(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[15]~q ),
	.av_readdata_pre_12(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[12]~q ),
	.av_readdata_pre_13(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[13]~q ),
	.av_readdata_pre_14(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[14]~q ),
	.clk(clk_clk));

first_nios2_system_altera_merlin_master_translator cpu_data_master_translator(
	.clr_break_line(clr_break_line),
	.reset(r_sync_rst),
	.d_read(d_read),
	.read_accepted1(\cpu_data_master_translator|read_accepted~q ),
	.uav_read(\cpu_data_master_translator|uav_read~0_combout ),
	.WideOr1(WideOr13),
	.WideOr0(\cmd_demux|WideOr0~3_combout ),
	.WideOr01(\cmd_demux|WideOr0~6_combout ),
	.av_waitrequest(cpu_data_master_waitrequest),
	.clk(clk_clk));

first_nios2_system_altera_merlin_slave_agent_13 rtd2_s1_agent(
	.mem_used_1(\rtd2_s1_agent_rsp_fifo|mem_used[1]~q ),
	.always1(\router|always1~12_combout ),
	.m0_write(\rtd2_s1_agent|m0_write~0_combout ));

first_nios2_system_altera_avalon_sc_fifo_12 rtd1_s1_agent_rsp_fifo(
	.reset(r_sync_rst),
	.read_latency_shift_reg_0(\rtd1_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_used_1(\rtd1_s1_agent_rsp_fifo|mem_used[1]~q ),
	.sink_ready(\cmd_demux|sink_ready~7_combout ),
	.sink_ready1(\cmd_demux|sink_ready~17_combout ),
	.clk(clk_clk));

first_nios2_system_altera_merlin_slave_agent_12 rtd1_s1_agent(
	.mem_used_1(\rtd1_s1_agent_rsp_fifo|mem_used[1]~q ),
	.always1(\router|always1~11_combout ),
	.m0_write(\rtd1_s1_agent|m0_write~0_combout ));

first_nios2_system_altera_avalon_sc_fifo_1 camdata2_s1_agent_rsp_fifo(
	.reset(r_sync_rst),
	.read_latency_shift_reg_0(\camdata2_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_used_1(\camdata2_s1_agent_rsp_fifo|mem_used[1]~q ),
	.sink_ready(\cmd_demux|sink_ready~6_combout ),
	.sink_ready1(\cmd_demux|sink_ready~16_combout ),
	.clk(clk_clk));

first_nios2_system_altera_merlin_slave_agent_1 camdata2_s1_agent(
	.always1(\router|always1~9_combout ),
	.mem_used_1(\camdata2_s1_agent_rsp_fifo|mem_used[1]~q ),
	.m0_write(\camdata2_s1_agent|m0_write~0_combout ));

first_nios2_system_altera_avalon_sc_fifo camdata1_s1_agent_rsp_fifo(
	.reset(r_sync_rst),
	.read_latency_shift_reg_0(\camdata1_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_used_1(\camdata1_s1_agent_rsp_fifo|mem_used[1]~q ),
	.sink_ready(\cmd_demux|sink_ready~0_combout ),
	.sink_ready1(\cmd_demux|sink_ready~12_combout ),
	.clk(clk_clk));

first_nios2_system_altera_merlin_slave_agent camdata1_s1_agent(
	.mem_used_1(\camdata1_s1_agent_rsp_fifo|mem_used[1]~q ),
	.always1(\router|always1~3_combout ),
	.m0_write(\camdata1_s1_agent|m0_write~0_combout ));

first_nios2_system_altera_avalon_sc_fifo_6 download2_s1_agent_rsp_fifo(
	.reset(r_sync_rst),
	.wait_latency_counter_1(\download2_s1_translator|wait_latency_counter[1]~q ),
	.mem_used_1(\download2_s1_agent_rsp_fifo|mem_used[1]~q ),
	.Equal14(\router|Equal14~0_combout ),
	.m0_write(\download2_s1_agent|m0_write~0_combout ),
	.write(write),
	.wait_latency_counter_0(wait_latency_counter_01),
	.Equal2(\router|Equal2~1_combout ),
	.m0_write1(\tenout2_s1_agent|m0_write~0_combout ),
	.read_latency_shift_reg(read_latency_shift_reg),
	.read_latency_shift_reg_0(\download2_s1_translator|read_latency_shift_reg[0]~q ),
	.clk(clk_clk));

first_nios2_system_altera_avalon_sc_fifo_3 camstate2_s1_agent_rsp_fifo(
	.reset(r_sync_rst),
	.read_latency_shift_reg_0(\camstate2_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_used_1(\camstate2_s1_agent_rsp_fifo|mem_used[1]~q ),
	.av_waitrequest_generated(\camstate2_s1_translator|av_waitrequest_generated~0_combout ),
	.sink_ready(\cmd_demux|sink_ready~4_combout ),
	.sink_ready1(\cmd_demux|sink_ready~11_combout ),
	.clk(clk_clk));

first_nios2_system_altera_merlin_slave_agent_3 camstate2_s1_agent(
	.always1(\router|always1~1_combout ),
	.mem_used_1(\camstate2_s1_agent_rsp_fifo|mem_used[1]~q ),
	.always11(\router|always1~6_combout ),
	.m0_write(\camstate2_s1_agent|m0_write~0_combout ));

first_nios2_system_altera_avalon_sc_fifo_2 camstate1_s1_agent_rsp_fifo(
	.reset(r_sync_rst),
	.read_latency_shift_reg_0(read_latency_shift_reg_0),
	.mem_used_1(\camstate1_s1_agent_rsp_fifo|mem_used[1]~q ),
	.av_waitrequest_generated(\camstate1_s1_translator|av_waitrequest_generated~0_combout ),
	.sink_ready(\cmd_demux|sink_ready~3_combout ),
	.sink_ready1(\cmd_demux|sink_ready~10_combout ),
	.clk(clk_clk));

first_nios2_system_altera_merlin_slave_agent_2 camstate1_s1_agent(
	.Equal6(\router|Equal6~0_combout ),
	.always1(\router|always1~1_combout ),
	.mem_used_1(\camstate1_s1_agent_rsp_fifo|mem_used[1]~q ),
	.m0_write(\camstate1_s1_agent|m0_write~0_combout ));

first_nios2_system_altera_avalon_sc_fifo_14 start_s1_agent_rsp_fifo(
	.A_mem_baddr_4(A_mem_baddr_4),
	.A_mem_baddr_7(A_mem_baddr_7),
	.A_mem_baddr_6(A_mem_baddr_6),
	.reset(r_sync_rst),
	.wait_latency_counter_1(wait_latency_counter_14),
	.Equal2(\router|Equal2~1_combout ),
	.mem_used_1(\start_s1_agent_rsp_fifo|mem_used[1]~q ),
	.m0_write(m0_write),
	.wait_latency_counter_0(wait_latency_counter_05),
	.m0_write1(\tenout2_s1_agent|m0_write~0_combout ),
	.read_latency_shift_reg(read_latency_shift_reg),
	.read_latency_shift_reg_0(\start_s1_translator|read_latency_shift_reg[0]~q ),
	.av_waitrequest_generated(\start_s1_translator|av_waitrequest_generated~0_combout ),
	.clk(clk_clk));

first_nios2_system_altera_merlin_slave_agent_14 start_s1_agent(
	.A_mem_baddr_4(A_mem_baddr_4),
	.A_mem_baddr_7(A_mem_baddr_7),
	.A_mem_baddr_6(A_mem_baddr_6),
	.Equal2(\router|Equal2~1_combout ),
	.mem_used_1(\start_s1_agent_rsp_fifo|mem_used[1]~q ),
	.m0_write(m0_write));

first_nios2_system_altera_avalon_sc_fifo_13 rtd2_s1_agent_rsp_fifo(
	.reset(r_sync_rst),
	.read_latency_shift_reg_0(\rtd2_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_used_1(\rtd2_s1_agent_rsp_fifo|mem_used[1]~q ),
	.sink_ready(\cmd_demux|sink_ready~8_combout ),
	.sink_ready1(\cmd_demux|sink_ready~18_combout ),
	.clk(clk_clk));

first_nios2_system_altera_merlin_slave_agent_18 tenout2_s1_agent(
	.clr_break_line(clr_break_line),
	.d_write(d_write),
	.m0_write(\tenout2_s1_agent|m0_write~0_combout ),
	.always1(\router|always1~5_combout ),
	.mem_used_1(\tenout2_s1_agent_rsp_fifo|mem_used[1]~q ),
	.m0_write1(\tenout2_s1_agent|m0_write~1_combout ));

first_nios2_system_altera_avalon_sc_fifo_17 tenout1_s1_agent_rsp_fifo(
	.reset(r_sync_rst),
	.read_latency_shift_reg_0(\tenout1_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_used_1(\tenout1_s1_agent_rsp_fifo|mem_used[1]~q ),
	.sink_ready(\cmd_demux|sink_ready~1_combout ),
	.sink_ready1(\cmd_demux|sink_ready~13_combout ),
	.clk(clk_clk));

first_nios2_system_altera_merlin_slave_agent_17 tenout1_s1_agent(
	.always1(\router|always1~4_combout ),
	.mem_used_1(\tenout1_s1_agent_rsp_fifo|mem_used[1]~q ),
	.m0_write(\tenout1_s1_agent|m0_write~0_combout ));

first_nios2_system_altera_avalon_sc_fifo_8 hex2_s1_agent_rsp_fifo(
	.A_mem_baddr_7(A_mem_baddr_7),
	.reset(r_sync_rst),
	.wait_latency_counter_1(wait_latency_counter_12),
	.mem_used_1(mem_used_12),
	.always1(always1),
	.wait_latency_counter_0(wait_latency_counter_03),
	.m0_write(\tenout2_s1_agent|m0_write~0_combout ),
	.read_latency_shift_reg(read_latency_shift_reg),
	.read_latency_shift_reg_0(\hex2_s1_translator|read_latency_shift_reg[0]~q ),
	.write(\hex2_s1_agent_rsp_fifo|write~0_combout ),
	.av_waitrequest_generated(\hex2_s1_translator|av_waitrequest_generated~0_combout ),
	.clk(clk_clk));

first_nios2_system_altera_merlin_slave_agent_8 hex2_s1_agent(
	.A_mem_baddr_7(A_mem_baddr_7),
	.mem_used_1(mem_used_12),
	.always1(always1),
	.m0_write(\hex2_s1_agent|m0_write~0_combout ));

first_nios2_system_altera_avalon_sc_fifo_7 hex1_s1_agent_rsp_fifo(
	.reset(r_sync_rst),
	.wait_latency_counter_1(wait_latency_counter_11),
	.mem_used_1(mem_used_11),
	.Equal6(Equal6),
	.wait_latency_counter_0(wait_latency_counter_02),
	.m0_write(\tenout2_s1_agent|m0_write~0_combout ),
	.read_latency_shift_reg(read_latency_shift_reg),
	.read_latency_shift_reg_0(\hex1_s1_translator|read_latency_shift_reg[0]~q ),
	.write(\hex1_s1_agent_rsp_fifo|write~0_combout ),
	.av_waitrequest_generated(\hex1_s1_translator|av_waitrequest_generated~0_combout ),
	.clk(clk_clk));

first_nios2_system_altera_merlin_slave_agent_7 hex1_s1_agent(
	.mem_used_1(mem_used_11),
	.Equal6(Equal6),
	.m0_write(\hex1_s1_agent|m0_write~0_combout ));

first_nios2_system_first_nios2_system_mm_interconnect_0_router_001 router_001(
	.ic_fill_tag_5(ic_fill_tag_5),
	.ic_fill_tag_4(ic_fill_tag_4),
	.ic_fill_tag_3(ic_fill_tag_3),
	.ic_fill_tag_2(ic_fill_tag_2),
	.ic_fill_tag_1(ic_fill_tag_1),
	.ic_fill_tag_0(ic_fill_tag_0),
	.Equal1(\router_001|Equal1~0_combout ));

first_nios2_system_first_nios2_system_mm_interconnect_0_router router(
	.A_mem_baddr_4(A_mem_baddr_4),
	.A_mem_baddr_5(A_mem_baddr_5),
	.A_mem_baddr_8(A_mem_baddr_8),
	.A_mem_baddr_16(A_mem_baddr_16),
	.A_mem_baddr_15(A_mem_baddr_15),
	.A_mem_baddr_14(A_mem_baddr_14),
	.A_mem_baddr_13(A_mem_baddr_13),
	.Equal1(Equal1),
	.A_mem_baddr_12(A_mem_baddr_12),
	.A_mem_baddr_11(A_mem_baddr_11),
	.A_mem_baddr_10(A_mem_baddr_10),
	.A_mem_baddr_9(A_mem_baddr_9),
	.Equal2(Equal2),
	.A_mem_baddr_7(A_mem_baddr_7),
	.A_mem_baddr_6(A_mem_baddr_6),
	.Equal15(Equal15),
	.A_mem_baddr_3(A_mem_baddr_3),
	.Equal14(\router|Equal14~0_combout ),
	.Equal6(\router|Equal6~0_combout ),
	.Equal61(Equal6),
	.always1(always1),
	.Equal16(Equal16),
	.Equal21(\router|Equal2~1_combout ),
	.uav_read(\cpu_data_master_translator|uav_read~0_combout ),
	.Equal22(Equal21),
	.always11(\router|always1~1_combout ),
	.always12(always11),
	.src_channel_2(\router|src_channel[2]~2_combout ),
	.src_channel_21(\router|src_channel[2]~3_combout ),
	.Equal11(\router|Equal1~1_combout ),
	.always13(\router|always1~3_combout ),
	.always14(\router|always1~4_combout ),
	.always15(\router|always1~5_combout ),
	.always16(\router|always1~6_combout ),
	.always17(\router|always1~7_combout ),
	.always18(\router|always1~9_combout ),
	.always19(\router|always1~11_combout ),
	.always110(\router|always1~12_combout ),
	.always111(\router|always1~13_combout ));

first_nios2_system_altera_avalon_sc_fifo_18 tenout2_s1_agent_rsp_fifo(
	.reset(r_sync_rst),
	.read_latency_shift_reg_0(\tenout2_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_used_1(\tenout2_s1_agent_rsp_fifo|mem_used[1]~q ),
	.sink_ready(\cmd_demux|sink_ready~2_combout ),
	.sink_ready1(\cmd_demux|sink_ready~14_combout ),
	.clk(clk_clk));

first_nios2_system_first_nios2_system_mm_interconnect_0_cmd_mux_002_1 cmd_mux_003(
	.A_st_data_0(A_st_data_0),
	.A_mem_baddr_4(A_mem_baddr_4),
	.A_mem_baddr_5(A_mem_baddr_5),
	.A_mem_baddr_8(A_mem_baddr_8),
	.A_mem_baddr_14(A_mem_baddr_14),
	.A_mem_baddr_13(A_mem_baddr_13),
	.A_mem_baddr_12(A_mem_baddr_12),
	.A_mem_baddr_11(A_mem_baddr_11),
	.A_mem_baddr_10(A_mem_baddr_10),
	.A_mem_baddr_9(A_mem_baddr_9),
	.A_mem_baddr_7(A_mem_baddr_7),
	.A_mem_baddr_6(A_mem_baddr_6),
	.clr_break_line(clr_break_line),
	.A_mem_baddr_3(A_mem_baddr_3),
	.A_mem_baddr_2(A_mem_baddr_2),
	.r_sync_rst(r_sync_rst),
	.A_st_data_1(A_st_data_1),
	.A_st_data_2(A_st_data_2),
	.A_st_data_3(A_st_data_3),
	.A_st_data_4(A_st_data_4),
	.A_st_data_5(A_st_data_5),
	.A_st_data_6(A_st_data_6),
	.A_st_data_7(A_st_data_7),
	.cp_valid(cp_valid),
	.saved_grant_0(saved_grant_0),
	.src_channel_2(\router|src_channel[2]~2_combout ),
	.src_channel_21(\router|src_channel[2]~3_combout ),
	.Equal1(\router|Equal1~1_combout ),
	.has_pending_responses(\cpu_instruction_master_limiter|has_pending_responses~q ),
	.i_read(i_read),
	.ic_fill_tag_3(ic_fill_tag_3),
	.ic_fill_tag_2(ic_fill_tag_2),
	.ic_fill_tag_1(ic_fill_tag_1),
	.ic_fill_tag_0(ic_fill_tag_0),
	.Equal11(\router_001|Equal1~0_combout ),
	.saved_grant_1(\cmd_mux_003|saved_grant[1]~q ),
	.last_dest_id_3(\cpu_instruction_master_limiter|last_dest_id[3]~q ),
	.WideOr11(WideOr15),
	.read_latency_shift_reg(\onchip_mem_s1_translator|read_latency_shift_reg~0_combout ),
	.src3_valid(\cmd_demux|src3_valid~0_combout ),
	.src1_valid(\cmd_demux_001|src1_valid~0_combout ),
	.ic_fill_ap_offset_0(ic_fill_ap_offset_0),
	.ic_fill_line_0(ic_fill_line_0),
	.ic_fill_ap_offset_2(ic_fill_ap_offset_2),
	.ic_fill_ap_offset_1(ic_fill_ap_offset_1),
	.ic_fill_line_5(ic_fill_line_5),
	.ic_fill_line_4(ic_fill_line_4),
	.ic_fill_line_3(ic_fill_line_3),
	.ic_fill_line_2(ic_fill_line_2),
	.ic_fill_line_1(ic_fill_line_1),
	.A_mem_byte_en_0(A_mem_byte_en_0),
	.src_payload(src_payload44),
	.src_data_38(src_data_381),
	.src_data_39(src_data_391),
	.src_data_40(src_data_401),
	.src_data_41(src_data_411),
	.src_data_42(src_data_421),
	.src_data_43(src_data_431),
	.src_data_44(src_data_441),
	.src_data_45(src_data_451),
	.src_data_46(src_data_461),
	.src_data_47(src_data_47),
	.src_data_48(src_data_48),
	.src_data_49(src_data_49),
	.src_data_50(src_data_50),
	.src_data_32(src_data_321),
	.A_st_data_16(A_st_data_16),
	.src_payload1(src_payload47),
	.src_payload2(src_payload48),
	.src_payload3(src_payload49),
	.src_payload4(src_payload50),
	.src_payload5(src_payload51),
	.src_payload6(src_payload52),
	.src_payload7(src_payload53),
	.A_st_data_22(A_st_data_22),
	.src_payload8(src_payload54),
	.A_mem_byte_en_2(A_mem_byte_en_2),
	.src_data_34(src_data_34),
	.A_st_data_23(A_st_data_23),
	.src_payload9(src_payload55),
	.A_st_data_24(A_st_data_24),
	.src_payload10(src_payload56),
	.A_mem_byte_en_3(A_mem_byte_en_3),
	.src_data_35(src_data_35),
	.A_st_data_25(A_st_data_25),
	.src_payload11(src_payload57),
	.A_st_data_31(A_st_data_31),
	.src_payload12(src_payload58),
	.A_st_data_21(A_st_data_21),
	.src_payload13(src_payload59),
	.A_st_data_11(A_st_data_11),
	.src_payload14(src_payload60),
	.A_mem_byte_en_1(A_mem_byte_en_1),
	.src_data_33(src_data_33),
	.A_st_data_28(A_st_data_28),
	.src_payload15(src_payload61),
	.A_st_data_10(A_st_data_10),
	.src_payload16(src_payload62),
	.A_st_data_27(A_st_data_27),
	.src_payload17(src_payload63),
	.A_st_data_8(A_st_data_8),
	.src_payload18(src_payload64),
	.A_st_data_9(A_st_data_9),
	.src_payload19(src_payload65),
	.A_st_data_26(A_st_data_26),
	.src_payload20(src_payload66),
	.A_st_data_20(A_st_data_20),
	.src_payload21(src_payload67),
	.A_st_data_19(A_st_data_19),
	.src_payload22(src_payload68),
	.A_st_data_17(A_st_data_17),
	.src_payload23(src_payload69),
	.A_st_data_30(A_st_data_30),
	.src_payload24(src_payload70),
	.A_st_data_18(A_st_data_18),
	.src_payload25(src_payload71),
	.src_payload26(src_payload72),
	.A_st_data_15(A_st_data_15),
	.src_payload27(src_payload73),
	.A_st_data_12(A_st_data_12),
	.src_payload28(src_payload74),
	.A_st_data_13(A_st_data_13),
	.src_payload29(src_payload75),
	.A_st_data_14(A_st_data_14),
	.src_payload30(src_payload76),
	.A_st_data_29(A_st_data_29),
	.src_payload31(src_payload77),
	.clk_clk(clk_clk));

first_nios2_system_first_nios2_system_mm_interconnect_0_cmd_mux_002 cmd_mux_002(
	.A_st_data_0(A_st_data_0),
	.A_mem_baddr_4(A_mem_baddr_4),
	.A_mem_baddr_5(A_mem_baddr_5),
	.A_mem_baddr_8(A_mem_baddr_8),
	.A_mem_baddr_10(A_mem_baddr_10),
	.A_mem_baddr_9(A_mem_baddr_9),
	.A_mem_baddr_7(A_mem_baddr_7),
	.A_mem_baddr_6(A_mem_baddr_6),
	.clr_break_line(clr_break_line),
	.A_mem_baddr_3(A_mem_baddr_3),
	.A_mem_baddr_2(A_mem_baddr_2),
	.r_sync_rst(r_sync_rst),
	.A_st_data_1(A_st_data_1),
	.A_st_data_2(A_st_data_2),
	.A_st_data_3(A_st_data_3),
	.A_st_data_4(A_st_data_4),
	.A_st_data_5(A_st_data_5),
	.A_st_data_6(A_st_data_6),
	.A_st_data_7(A_st_data_7),
	.cp_valid(cp_valid),
	.W_debug_mode(W_debug_mode),
	.src_channel_2(\router|src_channel[2]~2_combout ),
	.src_channel_21(\router|src_channel[2]~3_combout ),
	.Equal1(\router|Equal1~1_combout ),
	.saved_grant_0(saved_grant_01),
	.write(\cpu_debug_mem_slave_agent_rsp_fifo|write~0_combout ),
	.saved_grant_1(\cmd_mux_002|saved_grant[1]~q ),
	.last_dest_id_2(\cpu_instruction_master_limiter|last_dest_id[2]~q ),
	.has_pending_responses(\cpu_instruction_master_limiter|has_pending_responses~q ),
	.i_read(i_read),
	.Equal11(\router_001|Equal1~0_combout ),
	.WideOr11(WideOr14),
	.src2_valid(\cmd_demux|src2_valid~0_combout ),
	.src0_valid(\cmd_demux_001|src0_valid~0_combout ),
	.src_payload(src_payload),
	.ic_fill_ap_offset_0(ic_fill_ap_offset_0),
	.src_data_38(src_data_38),
	.ic_fill_line_0(ic_fill_line_0),
	.src_data_41(src_data_41),
	.ic_fill_ap_offset_2(ic_fill_ap_offset_2),
	.src_data_40(src_data_40),
	.ic_fill_ap_offset_1(ic_fill_ap_offset_1),
	.src_data_39(src_data_39),
	.ic_fill_line_5(ic_fill_line_5),
	.src_data_46(src_data_46),
	.ic_fill_line_4(ic_fill_line_4),
	.src_data_45(src_data_45),
	.ic_fill_line_3(ic_fill_line_3),
	.src_data_44(src_data_44),
	.ic_fill_line_2(ic_fill_line_2),
	.src_data_43(src_data_43),
	.ic_fill_line_1(ic_fill_line_1),
	.src_data_42(src_data_42),
	.src_payload1(src_payload1),
	.src_payload2(src_payload7),
	.A_mem_byte_en_0(A_mem_byte_en_0),
	.src_data_32(src_data_32),
	.src_payload3(src_payload45),
	.A_st_data_16(A_st_data_16),
	.src_payload4(src_payload46),
	.A_st_data_22(A_st_data_22),
	.A_mem_byte_en_2(A_mem_byte_en_2),
	.A_st_data_23(A_st_data_23),
	.A_st_data_24(A_st_data_24),
	.A_mem_byte_en_3(A_mem_byte_en_3),
	.A_st_data_25(A_st_data_25),
	.A_st_data_31(A_st_data_31),
	.A_st_data_21(A_st_data_21),
	.A_st_data_11(A_st_data_11),
	.A_mem_byte_en_1(A_mem_byte_en_1),
	.A_st_data_28(A_st_data_28),
	.A_st_data_10(A_st_data_10),
	.A_st_data_27(A_st_data_27),
	.A_st_data_8(A_st_data_8),
	.A_st_data_9(A_st_data_9),
	.A_st_data_26(A_st_data_26),
	.A_st_data_20(A_st_data_20),
	.A_st_data_19(A_st_data_19),
	.A_st_data_17(A_st_data_17),
	.A_st_data_30(A_st_data_30),
	.A_st_data_18(A_st_data_18),
	.A_st_data_15(A_st_data_15),
	.A_st_data_12(A_st_data_12),
	.A_st_data_13(A_st_data_13),
	.A_st_data_14(A_st_data_14),
	.A_st_data_29(A_st_data_29),
	.src_payload5(src_payload78),
	.src_payload6(src_payload79),
	.src_data_34(src_data_341),
	.src_payload7(src_payload80),
	.src_payload8(src_payload81),
	.src_payload9(src_payload82),
	.src_payload10(src_payload83),
	.src_payload11(src_payload84),
	.src_payload12(src_payload85),
	.src_payload13(src_payload86),
	.src_payload14(src_payload87),
	.src_payload15(src_payload88),
	.src_data_35(src_data_351),
	.src_payload16(src_payload89),
	.src_payload17(src_payload90),
	.src_payload18(src_payload91),
	.src_payload19(src_payload92),
	.src_payload20(src_payload93),
	.src_payload21(src_payload94),
	.src_payload22(src_payload95),
	.src_data_33(src_data_331),
	.src_payload23(src_payload96),
	.src_payload24(src_payload97),
	.src_payload25(src_payload98),
	.src_payload26(src_payload99),
	.src_payload27(src_payload100),
	.src_payload28(src_payload101),
	.src_payload29(src_payload102),
	.src_payload30(src_payload103),
	.src_payload31(src_payload104),
	.src_payload32(src_payload105),
	.clk_clk(clk_clk));

first_nios2_system_first_nios2_system_mm_interconnect_0_cmd_demux_001 cmd_demux_001(
	.clr_break_line(clr_break_line),
	.write(\cpu_debug_mem_slave_agent_rsp_fifo|write~0_combout ),
	.saved_grant_1(\cmd_mux_002|saved_grant[1]~q ),
	.last_dest_id_2(\cpu_instruction_master_limiter|last_dest_id[2]~q ),
	.has_pending_responses(\cpu_instruction_master_limiter|has_pending_responses~q ),
	.i_read(i_read),
	.Equal1(\router_001|Equal1~0_combout ),
	.saved_grant_11(\cmd_mux_003|saved_grant[1]~q ),
	.last_dest_id_3(\cpu_instruction_master_limiter|last_dest_id[3]~q ),
	.read_latency_shift_reg(\onchip_mem_s1_translator|read_latency_shift_reg~0_combout ),
	.src1_valid(\cmd_demux_001|src1_valid~0_combout ),
	.src0_valid(\cmd_demux_001|src0_valid~0_combout ),
	.WideOr0(WideOr0));

first_nios2_system_first_nios2_system_mm_interconnect_0_cmd_demux cmd_demux(
	.clr_break_line(clr_break_line),
	.wait_latency_counter_1(\download2_s1_translator|wait_latency_counter[1]~q ),
	.m0_write(\download2_s1_agent|m0_write~0_combout ),
	.wait_latency_counter_0(wait_latency_counter_01),
	.Equal6(\router|Equal6~0_combout ),
	.wait_latency_counter_11(wait_latency_counter_14),
	.m0_write1(m0_write),
	.wait_latency_counter_01(wait_latency_counter_05),
	.m0_write2(\tenout2_s1_agent|m0_write~0_combout ),
	.cp_valid(cp_valid),
	.write(\hex1_s1_agent_rsp_fifo|write~0_combout ),
	.write1(\hex2_s1_agent_rsp_fifo|write~0_combout ),
	.write2(\sys_clk_timer_s1_agent_rsp_fifo|write~0_combout ),
	.mem_used_1(mem_used_15),
	.saved_grant_0(saved_grant_0),
	.always1(\router|always1~1_combout ),
	.src_channel_2(\router|src_channel[2]~2_combout ),
	.src_channel_21(\router|src_channel[2]~3_combout ),
	.Equal1(\router|Equal1~1_combout ),
	.write3(\download1_s1_agent_rsp_fifo|write~1_combout ),
	.write4(\leds_s1_agent_rsp_fifo|write~0_combout ),
	.WideOr0(\cmd_demux|WideOr0~3_combout ),
	.mem_used_11(\camdata1_s1_agent_rsp_fifo|mem_used[1]~q ),
	.wait_latency_counter_12(\camdata1_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_02(\camdata1_s1_translator|wait_latency_counter[0]~q ),
	.always11(\router|always1~3_combout ),
	.sink_ready(\cmd_demux|sink_ready~0_combout ),
	.always12(\router|always1~4_combout ),
	.mem_used_12(\tenout1_s1_agent_rsp_fifo|mem_used[1]~q ),
	.wait_latency_counter_13(\tenout1_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_03(\tenout1_s1_translator|wait_latency_counter[0]~q ),
	.sink_ready1(\cmd_demux|sink_ready~1_combout ),
	.always13(\router|always1~5_combout ),
	.mem_used_13(\tenout2_s1_agent_rsp_fifo|mem_used[1]~q ),
	.wait_latency_counter_14(\tenout2_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_04(\tenout2_s1_translator|wait_latency_counter[0]~q ),
	.sink_ready2(\cmd_demux|sink_ready~2_combout ),
	.mem_used_14(\camstate1_s1_agent_rsp_fifo|mem_used[1]~q ),
	.av_waitrequest_generated(\camstate1_s1_translator|av_waitrequest_generated~0_combout ),
	.sink_ready3(\cmd_demux|sink_ready~3_combout ),
	.mem_used_15(\camstate2_s1_agent_rsp_fifo|mem_used[1]~q ),
	.always14(\router|always1~6_combout ),
	.av_waitrequest_generated1(\camstate2_s1_translator|av_waitrequest_generated~0_combout ),
	.sink_ready4(\cmd_demux|sink_ready~4_combout ),
	.av_waitrequest(av_waitrequest),
	.av_waitrequest1(av_waitrequest1),
	.mem_used_16(\sysid_control_slave_agent_rsp_fifo|mem_used[1]~q ),
	.wait_latency_counter_15(\sysid_control_slave_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_05(\sysid_control_slave_translator|wait_latency_counter[0]~q ),
	.always15(\router|always1~7_combout ),
	.sink_ready5(\cmd_demux|sink_ready~5_combout ),
	.always16(\router|always1~9_combout ),
	.mem_used_17(\camdata2_s1_agent_rsp_fifo|mem_used[1]~q ),
	.wait_latency_counter_16(\camdata2_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_06(\camdata2_s1_translator|wait_latency_counter[0]~q ),
	.sink_ready6(\cmd_demux|sink_ready~6_combout ),
	.mem_used_18(\rtd1_s1_agent_rsp_fifo|mem_used[1]~q ),
	.wait_latency_counter_17(\rtd1_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_07(\rtd1_s1_translator|wait_latency_counter[0]~q ),
	.always17(\router|always1~11_combout ),
	.sink_ready7(\cmd_demux|sink_ready~7_combout ),
	.mem_used_19(\rtd2_s1_agent_rsp_fifo|mem_used[1]~q ),
	.wait_latency_counter_18(\rtd2_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_08(\rtd2_s1_translator|wait_latency_counter[0]~q ),
	.always18(\router|always1~12_combout ),
	.sink_ready8(\cmd_demux|sink_ready~8_combout ),
	.saved_grant_01(saved_grant_01),
	.write5(\cpu_debug_mem_slave_agent_rsp_fifo|write~0_combout ),
	.WideOr01(\cmd_demux|WideOr0~6_combout ),
	.sink_ready9(\cmd_demux|sink_ready~10_combout ),
	.sink_ready10(\cmd_demux|sink_ready~11_combout ),
	.src3_valid(\cmd_demux|src3_valid~0_combout ),
	.sink_ready11(\cmd_demux|sink_ready~12_combout ),
	.sink_ready12(\cmd_demux|sink_ready~13_combout ),
	.sink_ready13(\cmd_demux|sink_ready~14_combout ),
	.sink_ready14(\cmd_demux|sink_ready~15_combout ),
	.sink_ready15(\cmd_demux|sink_ready~16_combout ),
	.sink_ready16(\cmd_demux|sink_ready~17_combout ),
	.sink_ready17(\cmd_demux|sink_ready~18_combout ),
	.src2_valid(\cmd_demux|src2_valid~0_combout ));

first_nios2_system_altera_merlin_traffic_limiter cpu_instruction_master_limiter(
	.clr_break_line(clr_break_line),
	.reset(r_sync_rst),
	.last_dest_id_2(\cpu_instruction_master_limiter|last_dest_id[2]~q ),
	.has_pending_responses1(\cpu_instruction_master_limiter|has_pending_responses~q ),
	.i_read(i_read),
	.cmd_sink_data({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\router_001|Equal1~0_combout ,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.last_dest_id_3(\cpu_instruction_master_limiter|last_dest_id[3]~q ),
	.save_dest_id(save_dest_id),
	.WideOr0(WideOr0),
	.nonposted_cmd_accepted1(nonposted_cmd_accepted),
	.src1_valid(\rsp_demux_002|src1_valid~0_combout ),
	.src1_valid1(\rsp_demux_003|src1_valid~0_combout ),
	.mem_61_0(\cpu_debug_mem_slave_agent_rsp_fifo|mem[0][61]~q ),
	.mem_61_01(\onchip_mem_s1_agent_rsp_fifo|mem[0][61]~q ),
	.suppress_change_dest_id(suppress_change_dest_id),
	.clk(clk_clk));

first_nios2_system_first_nios2_system_mm_interconnect_0_rsp_demux_002_1 rsp_demux_003(
	.read_latency_shift_reg_0(\onchip_mem_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_74_0(\onchip_mem_s1_agent_rsp_fifo|mem[0][74]~q ),
	.mem_56_0(\onchip_mem_s1_agent_rsp_fifo|mem[0][56]~q ),
	.src0_valid(src0_valid1),
	.src1_valid(\rsp_demux_003|src1_valid~0_combout ));

first_nios2_system_first_nios2_system_mm_interconnect_0_rsp_demux_002 rsp_demux_002(
	.read_latency_shift_reg_0(\cpu_debug_mem_slave_translator|read_latency_shift_reg[0]~q ),
	.mem_74_0(\cpu_debug_mem_slave_agent_rsp_fifo|mem[0][74]~q ),
	.mem_56_0(\cpu_debug_mem_slave_agent_rsp_fifo|mem[0][56]~q ),
	.src0_valid(src0_valid),
	.src1_valid(\rsp_demux_002|src1_valid~0_combout ));

first_nios2_system_first_nios2_system_mm_interconnect_0_rsp_mux_001 rsp_mux_001(
	.q_a_0(q_a_0),
	.q_a_1(q_a_1),
	.q_a_2(q_a_2),
	.q_a_3(q_a_3),
	.q_a_4(q_a_4),
	.q_a_5(q_a_5),
	.q_a_6(q_a_6),
	.q_a_7(q_a_7),
	.q_a_22(q_a_22),
	.q_a_23(q_a_23),
	.q_a_24(q_a_24),
	.q_a_25(q_a_25),
	.q_a_31(q_a_31),
	.q_a_21(q_a_21),
	.q_a_11(q_a_11),
	.q_a_28(q_a_28),
	.q_a_10(q_a_10),
	.q_a_27(q_a_27),
	.q_a_8(q_a_8),
	.q_a_9(q_a_9),
	.q_a_26(q_a_26),
	.q_a_20(q_a_20),
	.q_a_19(q_a_19),
	.q_a_17(q_a_17),
	.q_a_30(q_a_30),
	.q_a_18(q_a_18),
	.q_a_16(q_a_16),
	.q_a_15(q_a_15),
	.q_a_12(q_a_12),
	.q_a_13(q_a_13),
	.q_a_14(q_a_14),
	.q_a_29(q_a_29),
	.src1_valid(\rsp_demux_002|src1_valid~0_combout ),
	.src1_valid1(\rsp_demux_003|src1_valid~0_combout ),
	.av_readdata_pre_0(\cpu_debug_mem_slave_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_1(\cpu_debug_mem_slave_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_2(\cpu_debug_mem_slave_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_3(\cpu_debug_mem_slave_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_4(\cpu_debug_mem_slave_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_5(\cpu_debug_mem_slave_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_6(\cpu_debug_mem_slave_translator|av_readdata_pre[6]~q ),
	.av_readdata_pre_7(\cpu_debug_mem_slave_translator|av_readdata_pre[7]~q ),
	.av_readdata_pre_22(av_readdata_pre_221),
	.av_readdata_pre_23(av_readdata_pre_23),
	.av_readdata_pre_24(av_readdata_pre_24),
	.av_readdata_pre_25(av_readdata_pre_25),
	.av_readdata_pre_31(av_readdata_pre_31),
	.av_readdata_pre_21(av_readdata_pre_21),
	.av_readdata_pre_11(av_readdata_pre_11),
	.av_readdata_pre_28(av_readdata_pre_28),
	.av_readdata_pre_10(av_readdata_pre_10),
	.av_readdata_pre_27(av_readdata_pre_27),
	.av_readdata_pre_8(av_readdata_pre_8),
	.av_readdata_pre_9(av_readdata_pre_9),
	.av_readdata_pre_26(av_readdata_pre_26),
	.av_readdata_pre_20(av_readdata_pre_201),
	.av_readdata_pre_19(av_readdata_pre_191),
	.av_readdata_pre_17(av_readdata_pre_17),
	.av_readdata_pre_30(av_readdata_pre_30),
	.av_readdata_pre_18(av_readdata_pre_18),
	.av_readdata_pre_16(av_readdata_pre_16),
	.av_readdata_pre_15(av_readdata_pre_15),
	.av_readdata_pre_12(av_readdata_pre_12),
	.av_readdata_pre_13(av_readdata_pre_13),
	.av_readdata_pre_14(av_readdata_pre_14),
	.av_readdata_pre_29(av_readdata_pre_29),
	.WideOr11(WideOr16),
	.src_data_26(src_data_26),
	.src_data_25(src_data_25),
	.src_data_24(src_data_24),
	.src_data_23(src_data_23),
	.src_data_22(src_data_22),
	.src_data_1(src_data_11),
	.src_data_0(src_data_01),
	.src_data_2(src_data_21),
	.src_data_3(src_data_31),
	.src_data_4(src_data_4),
	.src_data_5(src_data_5),
	.src_data_28(src_data_28),
	.src_data_31(src_data_311),
	.src_data_27(src_data_27),
	.src_data_29(src_data_29),
	.src_data_30(src_data_30),
	.src_data_11(src_data_111),
	.src_data_12(src_data_12),
	.src_data_13(src_data_13),
	.src_data_14(src_data_14),
	.src_data_15(src_data_15),
	.src_data_16(src_data_16),
	.src_data_9(src_data_9),
	.src_data_21(src_data_211),
	.src_data_6(src_data_6),
	.src_data_8(src_data_8),
	.src_data_17(src_data_17),
	.src_data_18(src_data_18),
	.src_data_10(src_data_10),
	.src_data_7(src_data_7),
	.src_data_20(src_data_20),
	.src_data_19(src_data_19));

first_nios2_system_first_nios2_system_mm_interconnect_0_rsp_mux rsp_mux(
	.av_readdata_pre_0(\download1_s1_translator|av_readdata_pre[0]~q ),
	.q_a_0(q_a_0),
	.av_readdata_pre_01(\download2_s1_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_02(\hex1_s1_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_03(\hex2_s1_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_04(\start_s1_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_05(\leds_s1_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_06(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_1(\leds_s1_translator|av_readdata_pre[1]~q ),
	.q_a_1(q_a_1),
	.av_readdata_pre_11(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_12(\hex1_s1_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_13(\hex2_s1_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_2(\leds_s1_translator|av_readdata_pre[2]~q ),
	.q_a_2(q_a_2),
	.av_readdata_pre_21(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_22(\hex1_s1_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_23(\hex2_s1_translator|av_readdata_pre[2]~q ),
	.q_a_3(q_a_3),
	.av_readdata_pre_3(\hex2_s1_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_31(\leds_s1_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_32(\hex1_s1_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_33(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_4(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_41(\leds_s1_translator|av_readdata_pre[4]~q ),
	.q_a_4(q_a_4),
	.av_readdata_pre_42(\hex1_s1_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_43(\hex2_s1_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_5(\hex2_s1_translator|av_readdata_pre[5]~q ),
	.q_a_5(q_a_5),
	.av_readdata_pre_51(\leds_s1_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_52(\hex1_s1_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_53(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[5]~q ),
	.q_a_6(q_a_6),
	.av_readdata_pre_6(\hex2_s1_translator|av_readdata_pre[6]~q ),
	.av_readdata_pre_61(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[6]~q ),
	.av_readdata_pre_62(\leds_s1_translator|av_readdata_pre[6]~q ),
	.av_readdata_pre_63(\hex1_s1_translator|av_readdata_pre[6]~q ),
	.q_a_7(q_a_7),
	.av_readdata_pre_7(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[7]~q ),
	.av_readdata_pre_71(\leds_s1_translator|av_readdata_pre[7]~q ),
	.av_readdata_pre_221(av_readdata_pre_22),
	.q_a_22(q_a_22),
	.q_a_23(q_a_23),
	.q_a_24(q_a_24),
	.q_a_25(q_a_25),
	.q_a_31(q_a_31),
	.q_a_21(q_a_21),
	.av_readdata_pre_211(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[21]~q ),
	.q_a_11(q_a_11),
	.q_a_28(q_a_28),
	.q_a_10(q_a_10),
	.q_a_27(q_a_27),
	.q_a_8(q_a_8),
	.q_a_9(q_a_9),
	.q_a_26(q_a_26),
	.av_readdata_pre_20(av_readdata_pre_20),
	.q_a_20(q_a_20),
	.av_readdata_pre_19(av_readdata_pre_19),
	.q_a_19(q_a_19),
	.q_a_17(q_a_17),
	.av_readdata_pre_17(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[17]~q ),
	.q_a_30(q_a_30),
	.q_a_18(q_a_18),
	.av_readdata_pre_18(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[18]~q ),
	.q_a_16(q_a_16),
	.av_readdata_pre_16(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[16]~q ),
	.q_a_15(q_a_15),
	.q_a_12(q_a_12),
	.q_a_13(q_a_13),
	.q_a_14(q_a_14),
	.q_a_29(q_a_29),
	.read_latency_shift_reg_0(\download1_s1_translator|read_latency_shift_reg[0]~q ),
	.read_latency_shift_reg_01(read_latency_shift_reg_0),
	.read_latency_shift_reg_02(\camstate2_s1_translator|read_latency_shift_reg[0]~q ),
	.read_latency_shift_reg_03(\hex1_s1_translator|read_latency_shift_reg[0]~q ),
	.read_latency_shift_reg_04(\hex2_s1_translator|read_latency_shift_reg[0]~q ),
	.read_latency_shift_reg_05(\tenout1_s1_translator|read_latency_shift_reg[0]~q ),
	.read_latency_shift_reg_06(\tenout2_s1_translator|read_latency_shift_reg[0]~q ),
	.WideOr11(WideOr1),
	.read_latency_shift_reg_07(\camdata1_s1_translator|read_latency_shift_reg[0]~q ),
	.read_latency_shift_reg_08(\camdata2_s1_translator|read_latency_shift_reg[0]~q ),
	.read_latency_shift_reg_09(\rtd1_s1_translator|read_latency_shift_reg[0]~q ),
	.read_latency_shift_reg_010(\rtd2_s1_translator|read_latency_shift_reg[0]~q ),
	.read_latency_shift_reg_011(\start_s1_translator|read_latency_shift_reg[0]~q ),
	.WideOr12(WideOr11),
	.read_latency_shift_reg_012(\download2_s1_translator|read_latency_shift_reg[0]~q ),
	.src0_valid(src0_valid),
	.src0_valid1(src0_valid1),
	.read_latency_shift_reg_013(read_latency_shift_reg_01),
	.read_latency_shift_reg_014(\sysid_control_slave_translator|read_latency_shift_reg[0]~q ),
	.read_latency_shift_reg_015(\sys_clk_timer_s1_translator|read_latency_shift_reg[0]~q ),
	.read_latency_shift_reg_016(\leds_s1_translator|read_latency_shift_reg[0]~q ),
	.WideOr13(WideOr12),
	.WideOr14(WideOr13),
	.av_readdata_pre_07(\cpu_debug_mem_slave_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_08(\camstate2_s1_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_09(\tenout1_s1_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_010(\tenout2_s1_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_011(\camstate1_s1_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_012(\rtd2_s1_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_013(\rtd1_s1_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_014(\sys_clk_timer_s1_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_015(\camdata1_s1_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_016(\camdata2_s1_translator|av_readdata_pre[0]~q ),
	.src_data_0(src_data_0),
	.av_readdata_pre_14(\tenout2_s1_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_15(\cpu_debug_mem_slave_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_110(\camdata1_s1_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_111(\camstate2_s1_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_30(\sysid_control_slave_translator|av_readdata_pre[30]~q ),
	.src_payload(src_payload2),
	.av_readdata_pre_112(\sys_clk_timer_s1_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_113(\camdata2_s1_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_114(\camstate1_s1_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_115(\tenout1_s1_translator|av_readdata_pre[1]~q ),
	.src_data_1(src_data_1),
	.av_readdata_pre_24(\tenout2_s1_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_25(\cpu_debug_mem_slave_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_26(\camdata1_s1_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_27(\camstate2_s1_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_28(\sys_clk_timer_s1_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_29(\camdata2_s1_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_210(\camstate1_s1_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_212(\tenout1_s1_translator|av_readdata_pre[2]~q ),
	.src_data_2(src_data_2),
	.av_readdata_pre_34(\camdata2_s1_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_35(\tenout2_s1_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_36(\cpu_debug_mem_slave_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_37(\camdata1_s1_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_38(\tenout1_s1_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_39(\sys_clk_timer_s1_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_310(\camstate1_s1_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_311(\camstate2_s1_translator|av_readdata_pre[3]~q ),
	.src_data_3(src_data_3),
	.av_readdata_pre_44(\sys_clk_timer_s1_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_45(\cpu_debug_mem_slave_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_46(\camdata1_s1_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_47(\camdata2_s1_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_48(\camstate1_s1_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_49(\camstate2_s1_translator|av_readdata_pre[4]~q ),
	.src_payload1(src_payload3),
	.av_readdata_pre_54(\cpu_debug_mem_slave_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_55(\camdata1_s1_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_56(\camdata2_s1_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_57(\sys_clk_timer_s1_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_58(\camstate1_s1_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_59(\camstate2_s1_translator|av_readdata_pre[5]~q ),
	.src_payload2(src_payload4),
	.av_readdata_pre_64(\camdata1_s1_translator|av_readdata_pre[6]~q ),
	.av_readdata_pre_65(\sys_clk_timer_s1_translator|av_readdata_pre[6]~q ),
	.av_readdata_pre_66(\cpu_debug_mem_slave_translator|av_readdata_pre[6]~q ),
	.av_readdata_pre_67(\camdata2_s1_translator|av_readdata_pre[6]~q ),
	.src_payload3(src_payload5),
	.av_readdata_pre_72(\sys_clk_timer_s1_translator|av_readdata_pre[7]~q ),
	.av_readdata_pre_73(\cpu_debug_mem_slave_translator|av_readdata_pre[7]~q ),
	.src_payload4(src_payload6),
	.av_readdata_pre_222(av_readdata_pre_221),
	.src_payload5(src_payload8),
	.av_readdata_pre_231(av_readdata_pre_23),
	.src_payload6(src_payload9),
	.av_readdata_pre_241(av_readdata_pre_24),
	.src_payload7(src_payload10),
	.av_readdata_pre_251(av_readdata_pre_25),
	.src_payload8(src_payload11),
	.av_readdata_pre_312(av_readdata_pre_31),
	.src_payload9(src_payload12),
	.av_readdata_pre_213(av_readdata_pre_21),
	.src_payload10(src_payload13),
	.src_payload11(src_payload14),
	.av_readdata_pre_116(av_readdata_pre_11),
	.av_readdata_pre_117(\sys_clk_timer_s1_translator|av_readdata_pre[11]~q ),
	.src_payload12(src_payload15),
	.src_payload13(src_payload16),
	.av_readdata_pre_281(av_readdata_pre_28),
	.src_payload14(src_payload17),
	.av_readdata_pre_10(av_readdata_pre_10),
	.av_readdata_pre_101(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[10]~q ),
	.av_readdata_pre_102(\sys_clk_timer_s1_translator|av_readdata_pre[10]~q ),
	.src_payload15(src_payload18),
	.src_payload16(src_payload19),
	.av_readdata_pre_271(av_readdata_pre_27),
	.src_payload17(src_payload20),
	.av_readdata_pre_8(av_readdata_pre_8),
	.av_readdata_pre_81(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[8]~q ),
	.av_readdata_pre_82(\sys_clk_timer_s1_translator|av_readdata_pre[8]~q ),
	.src_payload18(src_payload21),
	.src_payload19(src_payload22),
	.av_readdata_pre_9(av_readdata_pre_9),
	.av_readdata_pre_91(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[9]~q ),
	.av_readdata_pre_92(\sys_clk_timer_s1_translator|av_readdata_pre[9]~q ),
	.src_payload20(src_payload23),
	.src_payload21(src_payload24),
	.av_readdata_pre_261(av_readdata_pre_26),
	.src_payload22(src_payload25),
	.av_readdata_pre_201(av_readdata_pre_201),
	.src_payload23(src_payload26),
	.av_readdata_pre_191(av_readdata_pre_191),
	.src_payload24(src_payload27),
	.av_readdata_pre_171(av_readdata_pre_17),
	.src_payload25(src_payload28),
	.src_payload26(src_payload29),
	.av_readdata_pre_301(av_readdata_pre_30),
	.src_payload27(src_payload30),
	.av_readdata_pre_181(av_readdata_pre_18),
	.src_payload28(src_payload31),
	.src_payload29(src_payload32),
	.av_readdata_pre_161(av_readdata_pre_16),
	.src_payload30(src_payload33),
	.src_payload31(src_payload34),
	.av_readdata_pre_151(av_readdata_pre_15),
	.av_readdata_pre_152(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[15]~q ),
	.av_readdata_pre_153(\sys_clk_timer_s1_translator|av_readdata_pre[15]~q ),
	.src_payload32(src_payload35),
	.src_payload33(src_payload36),
	.av_readdata_pre_121(av_readdata_pre_12),
	.av_readdata_pre_122(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[12]~q ),
	.av_readdata_pre_123(\sys_clk_timer_s1_translator|av_readdata_pre[12]~q ),
	.src_payload34(src_payload37),
	.src_payload35(src_payload38),
	.av_readdata_pre_131(av_readdata_pre_13),
	.av_readdata_pre_132(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[13]~q ),
	.av_readdata_pre_133(\sys_clk_timer_s1_translator|av_readdata_pre[13]~q ),
	.src_payload36(src_payload39),
	.src_payload37(src_payload40),
	.av_readdata_pre_141(av_readdata_pre_14),
	.av_readdata_pre_142(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[14]~q ),
	.av_readdata_pre_143(\sys_clk_timer_s1_translator|av_readdata_pre[14]~q ),
	.src_payload38(src_payload41),
	.src_payload39(src_payload42),
	.av_readdata_pre_291(av_readdata_pre_29),
	.src_payload40(src_payload43));

endmodule

module first_nios2_system_altera_avalon_sc_fifo (
	reset,
	read_latency_shift_reg_0,
	mem_used_1,
	sink_ready,
	sink_ready1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	read_latency_shift_reg_0;
output 	mem_used_1;
input 	sink_ready;
input 	sink_ready1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem_used[0]~1_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~0_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cyclonev_lcell_comb \mem_used[0]~1 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_1),
	.datac(!sink_ready),
	.datad(!\mem_used[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~1 .extended_lut = "off";
defparam \mem_used[0]~1 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \mem_used[0]~1 .shared_arith = "off";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cyclonev_lcell_comb \mem_used[1]~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_1),
	.datac(!sink_ready1),
	.datad(!\mem_used[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~0 .extended_lut = "off";
defparam \mem_used[1]~0 .lut_mask = 64'hAF3FAF3FAF3FAF3F;
defparam \mem_used[1]~0 .shared_arith = "off";

endmodule

module first_nios2_system_altera_avalon_sc_fifo_1 (
	reset,
	read_latency_shift_reg_0,
	mem_used_1,
	sink_ready,
	sink_ready1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	read_latency_shift_reg_0;
output 	mem_used_1;
input 	sink_ready;
input 	sink_ready1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem_used[0]~1_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~0_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cyclonev_lcell_comb \mem_used[0]~1 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_1),
	.datac(!sink_ready),
	.datad(!\mem_used[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~1 .extended_lut = "off";
defparam \mem_used[0]~1 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \mem_used[0]~1 .shared_arith = "off";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cyclonev_lcell_comb \mem_used[1]~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_1),
	.datac(!sink_ready1),
	.datad(!\mem_used[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~0 .extended_lut = "off";
defparam \mem_used[1]~0 .lut_mask = 64'hAF3FAF3FAF3FAF3F;
defparam \mem_used[1]~0 .shared_arith = "off";

endmodule

module first_nios2_system_altera_avalon_sc_fifo_2 (
	reset,
	read_latency_shift_reg_0,
	mem_used_1,
	av_waitrequest_generated,
	sink_ready,
	sink_ready1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	read_latency_shift_reg_0;
output 	mem_used_1;
input 	av_waitrequest_generated;
input 	sink_ready;
input 	sink_ready1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem_used[0]~1_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~0_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cyclonev_lcell_comb \mem_used[0]~1 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_1),
	.datac(!sink_ready1),
	.datad(!\mem_used[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~1 .extended_lut = "off";
defparam \mem_used[0]~1 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \mem_used[0]~1 .shared_arith = "off";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cyclonev_lcell_comb \mem_used[1]~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_1),
	.datac(!av_waitrequest_generated),
	.datad(!sink_ready),
	.datae(!\mem_used[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~0 .extended_lut = "off";
defparam \mem_used[1]~0 .lut_mask = 64'hAFFF3FFFAFFF3FFF;
defparam \mem_used[1]~0 .shared_arith = "off";

endmodule

module first_nios2_system_altera_avalon_sc_fifo_3 (
	reset,
	read_latency_shift_reg_0,
	mem_used_1,
	av_waitrequest_generated,
	sink_ready,
	sink_ready1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	read_latency_shift_reg_0;
output 	mem_used_1;
input 	av_waitrequest_generated;
input 	sink_ready;
input 	sink_ready1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem_used[0]~1_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~0_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cyclonev_lcell_comb \mem_used[0]~1 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_1),
	.datac(!sink_ready1),
	.datad(!\mem_used[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~1 .extended_lut = "off";
defparam \mem_used[0]~1 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \mem_used[0]~1 .shared_arith = "off";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cyclonev_lcell_comb \mem_used[1]~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_1),
	.datac(!av_waitrequest_generated),
	.datad(!sink_ready),
	.datae(!\mem_used[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~0 .extended_lut = "off";
defparam \mem_used[1]~0 .lut_mask = 64'hAFFF3FFFAFFF3FFF;
defparam \mem_used[1]~0 .shared_arith = "off";

endmodule

module first_nios2_system_altera_avalon_sc_fifo_4 (
	reset,
	uav_read,
	read_latency_shift_reg_0,
	mem_74_0,
	mem_56_0,
	saved_grant_0,
	waitrequest,
	mem_used_1,
	write,
	saved_grant_1,
	i_read,
	WideOr1,
	mem,
	mem_61_0,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	uav_read;
input 	read_latency_shift_reg_0;
output 	mem_74_0;
output 	mem_56_0;
input 	saved_grant_0;
input 	waitrequest;
output 	mem_used_1;
output 	write;
input 	saved_grant_1;
input 	i_read;
input 	WideOr1;
output 	mem;
output 	mem_61_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem[1][74]~q ;
wire \mem~1_combout ;
wire \mem_used[0]~2_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~0_combout ;
wire \mem[1][56]~q ;
wire \mem~2_combout ;
wire \mem_used[1]~1_combout ;
wire \mem[1][98]~q ;
wire \mem~3_combout ;


dffeas \mem[0][74] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~0_combout ),
	.q(mem_74_0),
	.prn(vcc));
defparam \mem[0][74] .is_wysiwyg = "true";
defparam \mem[0][74] .power_up = "low";

dffeas \mem[0][56] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~0_combout ),
	.q(mem_56_0),
	.prn(vcc));
defparam \mem[0][56] .is_wysiwyg = "true";
defparam \mem[0][56] .power_up = "low";

dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cyclonev_lcell_comb \write~0 (
	.dataa(!waitrequest),
	.datab(!mem_used_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write),
	.sumout(),
	.cout(),
	.shareout());
defparam \write~0 .extended_lut = "off";
defparam \write~0 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \write~0 .shared_arith = "off";

cyclonev_lcell_comb \mem~0 (
	.dataa(!uav_read),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!i_read),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(mem),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~0 .extended_lut = "off";
defparam \mem~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \mem~0 .shared_arith = "off";

dffeas \mem[0][61] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~0_combout ),
	.q(mem_61_0),
	.prn(vcc));
defparam \mem[0][61] .is_wysiwyg = "true";
defparam \mem[0][61] .power_up = "low";

dffeas \mem[1][74] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][74]~q ),
	.prn(vcc));
defparam \mem[1][74] .is_wysiwyg = "true";
defparam \mem[1][74] .power_up = "low";

cyclonev_lcell_comb \mem~1 (
	.dataa(!mem_used_1),
	.datab(!saved_grant_1),
	.datac(!\mem[1][74]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~1 .extended_lut = "off";
defparam \mem~1 .lut_mask = 64'h2727272727272727;
defparam \mem~1 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[0]~2 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!waitrequest),
	.datac(!mem_used_1),
	.datad(!WideOr1),
	.datae(!mem),
	.dataf(!\mem_used[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~2 .extended_lut = "off";
defparam \mem_used[0]~2 .lut_mask = 64'hFFACFFFFFFFFFFFF;
defparam \mem_used[0]~2 .shared_arith = "off";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cyclonev_lcell_comb \mem_used[1]~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!\mem_used[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~0 .extended_lut = "off";
defparam \mem_used[1]~0 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \mem_used[1]~0 .shared_arith = "off";

dffeas \mem[1][56] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][56]~q ),
	.prn(vcc));
defparam \mem[1][56] .is_wysiwyg = "true";
defparam \mem[1][56] .power_up = "low";

cyclonev_lcell_comb \mem~2 (
	.dataa(!mem_used_1),
	.datab(!mem),
	.datac(!\mem[1][56]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~2 .extended_lut = "off";
defparam \mem~2 .lut_mask = 64'h2727272727272727;
defparam \mem~2 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[1]~1 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!waitrequest),
	.datac(!mem_used_1),
	.datad(!WideOr1),
	.datae(!mem),
	.dataf(!\mem_used[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~1 .extended_lut = "off";
defparam \mem_used[1]~1 .lut_mask = 64'hFFAFFFFFFFCFFFFF;
defparam \mem_used[1]~1 .shared_arith = "off";

dffeas \mem[1][98] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][98]~q ),
	.prn(vcc));
defparam \mem[1][98] .is_wysiwyg = "true";
defparam \mem[1][98] .power_up = "low";

cyclonev_lcell_comb \mem~3 (
	.dataa(!saved_grant_0),
	.datab(!mem_used_1),
	.datac(!saved_grant_1),
	.datad(!\mem[1][98]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~3 .extended_lut = "off";
defparam \mem~3 .lut_mask = 64'h47FF47FF47FF47FF;
defparam \mem~3 .shared_arith = "off";

endmodule

module first_nios2_system_altera_avalon_sc_fifo_5 (
	mem_used_1,
	Equal15,
	wait_latency_counter_1,
	wait_latency_counter_0,
	reset,
	read_latency_shift_reg_0,
	m0_write,
	read_latency_shift_reg,
	write,
	read_latency_shift_reg1,
	clk)/* synthesis synthesis_greybox=1 */;
output 	mem_used_1;
input 	Equal15;
input 	wait_latency_counter_1;
input 	wait_latency_counter_0;
input 	reset;
input 	read_latency_shift_reg_0;
input 	m0_write;
input 	read_latency_shift_reg;
output 	write;
input 	read_latency_shift_reg1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \write~0_combout ;
wire \mem_used[0]~1_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~0_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cyclonev_lcell_comb \write~1 (
	.dataa(!wait_latency_counter_1),
	.datab(!wait_latency_counter_0),
	.datac(!mem_used_1),
	.datad(!Equal15),
	.datae(!m0_write),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write),
	.sumout(),
	.cout(),
	.shareout());
defparam \write~1 .extended_lut = "off";
defparam \write~1 .lut_mask = 64'hFBFFFEFFFBFFFEFF;
defparam \write~1 .shared_arith = "off";

cyclonev_lcell_comb \write~0 (
	.dataa(!wait_latency_counter_1),
	.datab(!wait_latency_counter_0),
	.datac(!mem_used_1),
	.datad(!Equal15),
	.datae(!m0_write),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\write~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \write~0 .extended_lut = "off";
defparam \write~0 .lut_mask = 64'hEBFFBEFFEBFFBEFF;
defparam \write~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[0]~1 (
	.dataa(!mem_used_1),
	.datab(!read_latency_shift_reg_0),
	.datac(!\mem_used[0]~q ),
	.datad(!read_latency_shift_reg1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~1 .extended_lut = "off";
defparam \mem_used[0]~1 .lut_mask = 64'hDFFFDFFFDFFFDFFF;
defparam \mem_used[0]~1 .shared_arith = "off";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cyclonev_lcell_comb \mem_used[1]~0 (
	.dataa(!mem_used_1),
	.datab(!read_latency_shift_reg_0),
	.datac(!\write~0_combout ),
	.datad(!\mem_used[0]~q ),
	.datae(!read_latency_shift_reg),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~0 .extended_lut = "off";
defparam \mem_used[1]~0 .lut_mask = 64'hCF5FFFFFCF5FFFFF;
defparam \mem_used[1]~0 .shared_arith = "off";

endmodule

module first_nios2_system_altera_avalon_sc_fifo_6 (
	reset,
	wait_latency_counter_1,
	mem_used_1,
	Equal14,
	m0_write,
	write,
	wait_latency_counter_0,
	Equal2,
	m0_write1,
	read_latency_shift_reg,
	read_latency_shift_reg_0,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	wait_latency_counter_1;
output 	mem_used_1;
input 	Equal14;
input 	m0_write;
output 	write;
input 	wait_latency_counter_0;
input 	Equal2;
input 	m0_write1;
input 	read_latency_shift_reg;
input 	read_latency_shift_reg_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \write~1_combout ;
wire \mem_used[0]~2_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~0_combout ;
wire \mem_used[1]~1_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cyclonev_lcell_comb \write~0 (
	.dataa(!wait_latency_counter_1),
	.datab(!m0_write),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write),
	.sumout(),
	.cout(),
	.shareout());
defparam \write~0 .extended_lut = "off";
defparam \write~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \write~0 .shared_arith = "off";

cyclonev_lcell_comb \write~1 (
	.dataa(!wait_latency_counter_0),
	.datab(!m0_write),
	.datac(!m0_write1),
	.datad(!read_latency_shift_reg),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\write~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \write~1 .extended_lut = "off";
defparam \write~1 .lut_mask = 64'h96FF96FF96FF96FF;
defparam \write~1 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[0]~2 (
	.dataa(!mem_used_1),
	.datab(!write),
	.datac(!read_latency_shift_reg_0),
	.datad(!\mem_used[0]~q ),
	.datae(!\write~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~2 .extended_lut = "off";
defparam \mem_used[0]~2 .lut_mask = 64'hF7FFFFFFF7FFFFFF;
defparam \mem_used[0]~2 .shared_arith = "off";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cyclonev_lcell_comb \mem_used[1]~0 (
	.dataa(!wait_latency_counter_1),
	.datab(!Equal2),
	.datac(!Equal14),
	.datad(!read_latency_shift_reg_0),
	.datae(!\mem_used[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~0 .extended_lut = "off";
defparam \mem_used[1]~0 .lut_mask = 64'hFFBFFFFFFFBFFFFF;
defparam \mem_used[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[1]~1 (
	.dataa(!mem_used_1),
	.datab(!read_latency_shift_reg_0),
	.datac(!\mem_used[0]~q ),
	.datad(!\write~1_combout ),
	.datae(!\mem_used[1]~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~1 .extended_lut = "off";
defparam \mem_used[1]~1 .lut_mask = 64'hFDFFFFFFFDFFFFFF;
defparam \mem_used[1]~1 .shared_arith = "off";

endmodule

module first_nios2_system_altera_avalon_sc_fifo_7 (
	reset,
	wait_latency_counter_1,
	mem_used_1,
	Equal6,
	wait_latency_counter_0,
	m0_write,
	read_latency_shift_reg,
	read_latency_shift_reg_0,
	write,
	av_waitrequest_generated,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	wait_latency_counter_1;
output 	mem_used_1;
input 	Equal6;
input 	wait_latency_counter_0;
input 	m0_write;
input 	read_latency_shift_reg;
input 	read_latency_shift_reg_0;
output 	write;
input 	av_waitrequest_generated;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem_used[0]~1_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~0_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cyclonev_lcell_comb \write~0 (
	.dataa(!wait_latency_counter_0),
	.datab(!wait_latency_counter_1),
	.datac(!mem_used_1),
	.datad(!Equal6),
	.datae(!m0_write),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write),
	.sumout(),
	.cout(),
	.shareout());
defparam \write~0 .extended_lut = "off";
defparam \write~0 .lut_mask = 64'hFDFFFEFFFDFFFEFF;
defparam \write~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[0]~1 (
	.dataa(!mem_used_1),
	.datab(!read_latency_shift_reg_0),
	.datac(!write),
	.datad(!read_latency_shift_reg),
	.datae(!\mem_used[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~1 .extended_lut = "off";
defparam \mem_used[0]~1 .lut_mask = 64'hDFFFFFFFDFFFFFFF;
defparam \mem_used[0]~1 .shared_arith = "off";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cyclonev_lcell_comb \mem_used[1]~0 (
	.dataa(!mem_used_1),
	.datab(!Equal6),
	.datac(!read_latency_shift_reg_0),
	.datad(!read_latency_shift_reg),
	.datae(!av_waitrequest_generated),
	.dataf(!\mem_used[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~0 .extended_lut = "off";
defparam \mem_used[1]~0 .lut_mask = 64'hF3FFFFFF77FFFFFF;
defparam \mem_used[1]~0 .shared_arith = "off";

endmodule

module first_nios2_system_altera_avalon_sc_fifo_8 (
	A_mem_baddr_7,
	reset,
	wait_latency_counter_1,
	mem_used_1,
	always1,
	wait_latency_counter_0,
	m0_write,
	read_latency_shift_reg,
	read_latency_shift_reg_0,
	write,
	av_waitrequest_generated,
	clk)/* synthesis synthesis_greybox=1 */;
input 	A_mem_baddr_7;
input 	reset;
input 	wait_latency_counter_1;
output 	mem_used_1;
input 	always1;
input 	wait_latency_counter_0;
input 	m0_write;
input 	read_latency_shift_reg;
input 	read_latency_shift_reg_0;
output 	write;
input 	av_waitrequest_generated;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem_used[0]~3_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~0_combout ;
wire \mem_used[1]~1_combout ;
wire \mem_used[1]~2_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cyclonev_lcell_comb \write~0 (
	.dataa(!A_mem_baddr_7),
	.datab(!wait_latency_counter_0),
	.datac(!wait_latency_counter_1),
	.datad(!mem_used_1),
	.datae(!always1),
	.dataf(!m0_write),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write),
	.sumout(),
	.cout(),
	.shareout());
defparam \write~0 .extended_lut = "off";
defparam \write~0 .lut_mask = 64'hFFFBFFFFFFFEFFFF;
defparam \write~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[0]~3 (
	.dataa(!mem_used_1),
	.datab(!read_latency_shift_reg_0),
	.datac(!write),
	.datad(!read_latency_shift_reg),
	.datae(!\mem_used[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~3 .extended_lut = "off";
defparam \mem_used[0]~3 .lut_mask = 64'hDFFFFFFFDFFFFFFF;
defparam \mem_used[0]~3 .shared_arith = "off";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cyclonev_lcell_comb \mem_used[1]~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!read_latency_shift_reg),
	.datac(!\mem_used[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~0 .extended_lut = "off";
defparam \mem_used[1]~0 .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \mem_used[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[1]~1 (
	.dataa(!A_mem_baddr_7),
	.datab(!wait_latency_counter_1),
	.datac(!always1),
	.datad(!av_waitrequest_generated),
	.datae(!\mem_used[1]~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~1 .extended_lut = "off";
defparam \mem_used[1]~1 .lut_mask = 64'hEFFFFFFFEFFFFFFF;
defparam \mem_used[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[1]~2 (
	.dataa(!mem_used_1),
	.datab(!read_latency_shift_reg_0),
	.datac(!\mem_used[0]~q ),
	.datad(!\mem_used[1]~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~2 .extended_lut = "off";
defparam \mem_used[1]~2 .lut_mask = 64'hFDFFFDFFFDFFFDFF;
defparam \mem_used[1]~2 .shared_arith = "off";

endmodule

module first_nios2_system_altera_avalon_sc_fifo_9 (
	A_mem_baddr_4,
	A_mem_baddr_3,
	reset,
	read_latency_shift_reg,
	read_latency_shift_reg_0,
	av_waitrequest,
	mem_used_1,
	always1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	A_mem_baddr_4;
input 	A_mem_baddr_3;
input 	reset;
input 	read_latency_shift_reg;
input 	read_latency_shift_reg_0;
input 	av_waitrequest;
output 	mem_used_1;
input 	always1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \write~0_combout ;
wire \mem_used[0]~1_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~0_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cyclonev_lcell_comb \write~0 (
	.dataa(!A_mem_baddr_3),
	.datab(!A_mem_baddr_4),
	.datac(!av_waitrequest),
	.datad(!always1),
	.datae(!read_latency_shift_reg),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\write~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \write~0 .extended_lut = "off";
defparam \write~0 .lut_mask = 64'hDFFFFFFFDFFFFFFF;
defparam \write~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[0]~1 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_1),
	.datac(!\mem_used[0]~q ),
	.datad(!\write~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~1 .extended_lut = "off";
defparam \mem_used[0]~1 .lut_mask = 64'h8BFF8BFF8BFF8BFF;
defparam \mem_used[0]~1 .shared_arith = "off";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cyclonev_lcell_comb \mem_used[1]~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_1),
	.datac(!\mem_used[0]~q ),
	.datad(!\write~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~0 .extended_lut = "off";
defparam \mem_used[1]~0 .lut_mask = 64'hA3FFA3FFA3FFA3FF;
defparam \mem_used[1]~0 .shared_arith = "off";

endmodule

module first_nios2_system_altera_avalon_sc_fifo_10 (
	reset,
	wait_latency_counter_1,
	mem_used_1,
	Equal16,
	wait_latency_counter_0,
	m0_write,
	read_latency_shift_reg,
	read_latency_shift_reg_0,
	write,
	av_waitrequest_generated,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	wait_latency_counter_1;
output 	mem_used_1;
input 	Equal16;
input 	wait_latency_counter_0;
input 	m0_write;
input 	read_latency_shift_reg;
input 	read_latency_shift_reg_0;
output 	write;
input 	av_waitrequest_generated;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem_used[0]~1_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~0_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cyclonev_lcell_comb \write~0 (
	.dataa(!wait_latency_counter_0),
	.datab(!wait_latency_counter_1),
	.datac(!mem_used_1),
	.datad(!Equal16),
	.datae(!m0_write),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write),
	.sumout(),
	.cout(),
	.shareout());
defparam \write~0 .extended_lut = "off";
defparam \write~0 .lut_mask = 64'hFDFFFEFFFDFFFEFF;
defparam \write~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[0]~1 (
	.dataa(!mem_used_1),
	.datab(!read_latency_shift_reg_0),
	.datac(!write),
	.datad(!read_latency_shift_reg),
	.datae(!\mem_used[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~1 .extended_lut = "off";
defparam \mem_used[0]~1 .lut_mask = 64'hDFFFFFFFDFFFFFFF;
defparam \mem_used[0]~1 .shared_arith = "off";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cyclonev_lcell_comb \mem_used[1]~0 (
	.dataa(!mem_used_1),
	.datab(!Equal16),
	.datac(!read_latency_shift_reg_0),
	.datad(!read_latency_shift_reg),
	.datae(!av_waitrequest_generated),
	.dataf(!\mem_used[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~0 .extended_lut = "off";
defparam \mem_used[1]~0 .lut_mask = 64'hF3FFFFFF77FFFFFF;
defparam \mem_used[1]~0 .shared_arith = "off";

endmodule

module first_nios2_system_altera_avalon_sc_fifo_11 (
	clr_break_line,
	reset,
	uav_read,
	read_latency_shift_reg_0,
	mem_74_0,
	mem_56_0,
	mem_used_1,
	saved_grant_0,
	i_read,
	saved_grant_1,
	WideOr1,
	mem,
	mem_61_0,
	clk)/* synthesis synthesis_greybox=1 */;
input 	clr_break_line;
input 	reset;
input 	uav_read;
input 	read_latency_shift_reg_0;
output 	mem_74_0;
output 	mem_56_0;
output 	mem_used_1;
input 	saved_grant_0;
input 	i_read;
input 	saved_grant_1;
input 	WideOr1;
output 	mem;
output 	mem_61_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem[1][74]~q ;
wire \mem~1_combout ;
wire \mem_used[0]~2_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~0_combout ;
wire \mem[1][56]~q ;
wire \mem~2_combout ;
wire \mem_used[1]~1_combout ;
wire \mem[1][98]~q ;
wire \mem~3_combout ;


dffeas \mem[0][74] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~0_combout ),
	.q(mem_74_0),
	.prn(vcc));
defparam \mem[0][74] .is_wysiwyg = "true";
defparam \mem[0][74] .power_up = "low";

dffeas \mem[0][56] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~0_combout ),
	.q(mem_56_0),
	.prn(vcc));
defparam \mem[0][56] .is_wysiwyg = "true";
defparam \mem[0][56] .power_up = "low";

dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cyclonev_lcell_comb \mem~0 (
	.dataa(!uav_read),
	.datab(!saved_grant_0),
	.datac(!i_read),
	.datad(!saved_grant_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(mem),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~0 .extended_lut = "off";
defparam \mem~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \mem~0 .shared_arith = "off";

dffeas \mem[0][61] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~0_combout ),
	.q(mem_61_0),
	.prn(vcc));
defparam \mem[0][61] .is_wysiwyg = "true";
defparam \mem[0][61] .power_up = "low";

dffeas \mem[1][74] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][74]~q ),
	.prn(vcc));
defparam \mem[1][74] .is_wysiwyg = "true";
defparam \mem[1][74] .power_up = "low";

cyclonev_lcell_comb \mem~1 (
	.dataa(!mem_used_1),
	.datab(!saved_grant_1),
	.datac(!\mem[1][74]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~1 .extended_lut = "off";
defparam \mem~1 .lut_mask = 64'h2727272727272727;
defparam \mem~1 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[0]~2 (
	.dataa(!clr_break_line),
	.datab(!read_latency_shift_reg_0),
	.datac(!mem_used_1),
	.datad(!WideOr1),
	.datae(!mem),
	.dataf(!\mem_used[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~2 .extended_lut = "off";
defparam \mem_used[0]~2 .lut_mask = 64'hDFD5FFFFFFFFFFFF;
defparam \mem_used[0]~2 .shared_arith = "off";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cyclonev_lcell_comb \mem_used[1]~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!\mem_used[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~0 .extended_lut = "off";
defparam \mem_used[1]~0 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \mem_used[1]~0 .shared_arith = "off";

dffeas \mem[1][56] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][56]~q ),
	.prn(vcc));
defparam \mem[1][56] .is_wysiwyg = "true";
defparam \mem[1][56] .power_up = "low";

cyclonev_lcell_comb \mem~2 (
	.dataa(!mem_used_1),
	.datab(!mem),
	.datac(!\mem[1][56]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~2 .extended_lut = "off";
defparam \mem~2 .lut_mask = 64'h2727272727272727;
defparam \mem~2 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[1]~1 (
	.dataa(!clr_break_line),
	.datab(!read_latency_shift_reg_0),
	.datac(!mem_used_1),
	.datad(!WideOr1),
	.datae(!mem),
	.dataf(!\mem_used[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~1 .extended_lut = "off";
defparam \mem_used[1]~1 .lut_mask = 64'hDFDFFFFFFF5FFFFF;
defparam \mem_used[1]~1 .shared_arith = "off";

dffeas \mem[1][98] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][98]~q ),
	.prn(vcc));
defparam \mem[1][98] .is_wysiwyg = "true";
defparam \mem[1][98] .power_up = "low";

cyclonev_lcell_comb \mem~3 (
	.dataa(!mem_used_1),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!\mem[1][98]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~3 .extended_lut = "off";
defparam \mem~3 .lut_mask = 64'h27FF27FF27FF27FF;
defparam \mem~3 .shared_arith = "off";

endmodule

module first_nios2_system_altera_avalon_sc_fifo_12 (
	reset,
	read_latency_shift_reg_0,
	mem_used_1,
	sink_ready,
	sink_ready1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	read_latency_shift_reg_0;
output 	mem_used_1;
input 	sink_ready;
input 	sink_ready1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem_used[0]~1_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~0_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cyclonev_lcell_comb \mem_used[0]~1 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_1),
	.datac(!sink_ready),
	.datad(!\mem_used[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~1 .extended_lut = "off";
defparam \mem_used[0]~1 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \mem_used[0]~1 .shared_arith = "off";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cyclonev_lcell_comb \mem_used[1]~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_1),
	.datac(!sink_ready1),
	.datad(!\mem_used[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~0 .extended_lut = "off";
defparam \mem_used[1]~0 .lut_mask = 64'hAF3FAF3FAF3FAF3F;
defparam \mem_used[1]~0 .shared_arith = "off";

endmodule

module first_nios2_system_altera_avalon_sc_fifo_13 (
	reset,
	read_latency_shift_reg_0,
	mem_used_1,
	sink_ready,
	sink_ready1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	read_latency_shift_reg_0;
output 	mem_used_1;
input 	sink_ready;
input 	sink_ready1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem_used[0]~1_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~0_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cyclonev_lcell_comb \mem_used[0]~1 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_1),
	.datac(!sink_ready),
	.datad(!\mem_used[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~1 .extended_lut = "off";
defparam \mem_used[0]~1 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \mem_used[0]~1 .shared_arith = "off";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cyclonev_lcell_comb \mem_used[1]~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_1),
	.datac(!sink_ready1),
	.datad(!\mem_used[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~0 .extended_lut = "off";
defparam \mem_used[1]~0 .lut_mask = 64'hAF3FAF3FAF3FAF3F;
defparam \mem_used[1]~0 .shared_arith = "off";

endmodule

module first_nios2_system_altera_avalon_sc_fifo_14 (
	A_mem_baddr_4,
	A_mem_baddr_7,
	A_mem_baddr_6,
	reset,
	wait_latency_counter_1,
	Equal2,
	mem_used_1,
	m0_write,
	wait_latency_counter_0,
	m0_write1,
	read_latency_shift_reg,
	read_latency_shift_reg_0,
	av_waitrequest_generated,
	clk)/* synthesis synthesis_greybox=1 */;
input 	A_mem_baddr_4;
input 	A_mem_baddr_7;
input 	A_mem_baddr_6;
input 	reset;
input 	wait_latency_counter_1;
input 	Equal2;
output 	mem_used_1;
input 	m0_write;
input 	wait_latency_counter_0;
input 	m0_write1;
input 	read_latency_shift_reg;
input 	read_latency_shift_reg_0;
input 	av_waitrequest_generated;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \write~0_combout ;
wire \mem_used[0]~3_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~0_combout ;
wire \mem_used[1]~1_combout ;
wire \mem_used[1]~2_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cyclonev_lcell_comb \write~0 (
	.dataa(!wait_latency_counter_0),
	.datab(!wait_latency_counter_1),
	.datac(!m0_write),
	.datad(!m0_write1),
	.datae(!read_latency_shift_reg),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\write~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \write~0 .extended_lut = "off";
defparam \write~0 .lut_mask = 64'hDFEFFFFFDFEFFFFF;
defparam \write~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[0]~3 (
	.dataa(!mem_used_1),
	.datab(!read_latency_shift_reg_0),
	.datac(!\mem_used[0]~q ),
	.datad(!\write~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~3 .extended_lut = "off";
defparam \mem_used[0]~3 .lut_mask = 64'hDFFFDFFFDFFFDFFF;
defparam \mem_used[0]~3 .shared_arith = "off";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cyclonev_lcell_comb \mem_used[1]~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!read_latency_shift_reg),
	.datac(!\mem_used[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~0 .extended_lut = "off";
defparam \mem_used[1]~0 .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \mem_used[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[1]~1 (
	.dataa(!A_mem_baddr_4),
	.datab(!A_mem_baddr_7),
	.datac(!A_mem_baddr_6),
	.datad(!Equal2),
	.datae(!\mem_used[1]~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~1 .extended_lut = "off";
defparam \mem_used[1]~1 .lut_mask = 64'hFBFFFFFFFBFFFFFF;
defparam \mem_used[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[1]~2 (
	.dataa(!mem_used_1),
	.datab(!read_latency_shift_reg_0),
	.datac(!av_waitrequest_generated),
	.datad(!\mem_used[0]~q ),
	.datae(!\mem_used[1]~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~2 .extended_lut = "off";
defparam \mem_used[1]~2 .lut_mask = 64'hFFDFFFFFFFDFFFFF;
defparam \mem_used[1]~2 .shared_arith = "off";

endmodule

module first_nios2_system_altera_avalon_sc_fifo_15 (
	reset,
	m0_write,
	read_latency_shift_reg,
	read_latency_shift_reg_0,
	Equal2,
	wait_latency_counter_0,
	mem_used_1,
	wait_latency_counter_1,
	write,
	av_waitrequest_generated,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	m0_write;
input 	read_latency_shift_reg;
input 	read_latency_shift_reg_0;
input 	Equal2;
input 	wait_latency_counter_0;
output 	mem_used_1;
input 	wait_latency_counter_1;
output 	write;
input 	av_waitrequest_generated;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem_used[0]~1_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~0_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cyclonev_lcell_comb \write~0 (
	.dataa(!m0_write),
	.datab(!Equal2),
	.datac(!wait_latency_counter_0),
	.datad(!mem_used_1),
	.datae(!wait_latency_counter_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write),
	.sumout(),
	.cout(),
	.shareout());
defparam \write~0 .extended_lut = "off";
defparam \write~0 .lut_mask = 64'hFFFFFF7BFFFFFF7B;
defparam \write~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[0]~1 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_1),
	.datac(!write),
	.datad(!read_latency_shift_reg),
	.datae(!\mem_used[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~1 .extended_lut = "off";
defparam \mem_used[0]~1 .lut_mask = 64'hBFFFFFFFBFFFFFFF;
defparam \mem_used[0]~1 .shared_arith = "off";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cyclonev_lcell_comb \mem_used[1]~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!Equal2),
	.datac(!mem_used_1),
	.datad(!read_latency_shift_reg),
	.datae(!av_waitrequest_generated),
	.dataf(!\mem_used[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~0 .extended_lut = "off";
defparam \mem_used[1]~0 .lut_mask = 64'hAFFFFFFF3FFFFFFF;
defparam \mem_used[1]~0 .shared_arith = "off";

endmodule

module first_nios2_system_altera_avalon_sc_fifo_16 (
	reset,
	read_latency_shift_reg_0,
	mem_used_1,
	sink_ready,
	sink_ready1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	read_latency_shift_reg_0;
output 	mem_used_1;
input 	sink_ready;
input 	sink_ready1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem_used[0]~1_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~0_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cyclonev_lcell_comb \mem_used[0]~1 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_1),
	.datac(!sink_ready),
	.datad(!\mem_used[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~1 .extended_lut = "off";
defparam \mem_used[0]~1 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \mem_used[0]~1 .shared_arith = "off";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cyclonev_lcell_comb \mem_used[1]~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_1),
	.datac(!sink_ready1),
	.datad(!\mem_used[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~0 .extended_lut = "off";
defparam \mem_used[1]~0 .lut_mask = 64'hAF3FAF3FAF3FAF3F;
defparam \mem_used[1]~0 .shared_arith = "off";

endmodule

module first_nios2_system_altera_avalon_sc_fifo_17 (
	reset,
	read_latency_shift_reg_0,
	mem_used_1,
	sink_ready,
	sink_ready1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	read_latency_shift_reg_0;
output 	mem_used_1;
input 	sink_ready;
input 	sink_ready1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem_used[0]~1_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~0_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cyclonev_lcell_comb \mem_used[0]~1 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_1),
	.datac(!sink_ready),
	.datad(!\mem_used[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~1 .extended_lut = "off";
defparam \mem_used[0]~1 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \mem_used[0]~1 .shared_arith = "off";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cyclonev_lcell_comb \mem_used[1]~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_1),
	.datac(!sink_ready1),
	.datad(!\mem_used[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~0 .extended_lut = "off";
defparam \mem_used[1]~0 .lut_mask = 64'hAF3FAF3FAF3FAF3F;
defparam \mem_used[1]~0 .shared_arith = "off";

endmodule

module first_nios2_system_altera_avalon_sc_fifo_18 (
	reset,
	read_latency_shift_reg_0,
	mem_used_1,
	sink_ready,
	sink_ready1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	read_latency_shift_reg_0;
output 	mem_used_1;
input 	sink_ready;
input 	sink_ready1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem_used[0]~1_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~0_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cyclonev_lcell_comb \mem_used[0]~1 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_1),
	.datac(!sink_ready),
	.datad(!\mem_used[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~1 .extended_lut = "off";
defparam \mem_used[0]~1 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \mem_used[0]~1 .shared_arith = "off";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cyclonev_lcell_comb \mem_used[1]~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_1),
	.datac(!sink_ready1),
	.datad(!\mem_used[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~0 .extended_lut = "off";
defparam \mem_used[1]~0 .lut_mask = 64'hAF3FAF3FAF3FAF3F;
defparam \mem_used[1]~0 .shared_arith = "off";

endmodule

module first_nios2_system_altera_merlin_master_agent (
	clr_break_line,
	d_write,
	d_read,
	read_accepted,
	cp_valid)/* synthesis synthesis_greybox=1 */;
input 	clr_break_line;
input 	d_write;
input 	d_read;
input 	read_accepted;
output 	cp_valid;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \cp_valid~0 (
	.dataa(!clr_break_line),
	.datab(!d_write),
	.datac(!d_read),
	.datad(!read_accepted),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cp_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_valid~0 .extended_lut = "off";
defparam \cp_valid~0 .lut_mask = 64'hFF7FFF7FFF7FFF7F;
defparam \cp_valid~0 .shared_arith = "off";

endmodule

module first_nios2_system_altera_merlin_master_translator (
	clr_break_line,
	reset,
	d_read,
	read_accepted1,
	uav_read,
	WideOr1,
	WideOr0,
	WideOr01,
	av_waitrequest,
	clk)/* synthesis synthesis_greybox=1 */;
input 	clr_break_line;
input 	reset;
input 	d_read;
output 	read_accepted1;
output 	uav_read;
input 	WideOr1;
input 	WideOr0;
input 	WideOr01;
output 	av_waitrequest;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read_accepted~0_combout ;


dffeas read_accepted(
	.clk(clk),
	.d(\read_accepted~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_accepted1),
	.prn(vcc));
defparam read_accepted.is_wysiwyg = "true";
defparam read_accepted.power_up = "low";

cyclonev_lcell_comb \uav_read~0 (
	.dataa(!d_read),
	.datab(!read_accepted1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(uav_read),
	.sumout(),
	.cout(),
	.shareout());
defparam \uav_read~0 .extended_lut = "off";
defparam \uav_read~0 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \uav_read~0 .shared_arith = "off";

cyclonev_lcell_comb \av_waitrequest~0 (
	.dataa(!clr_break_line),
	.datab(!d_read),
	.datac(!WideOr1),
	.datad(!WideOr0),
	.datae(!WideOr01),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(av_waitrequest),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_waitrequest~0 .extended_lut = "off";
defparam \av_waitrequest~0 .lut_mask = 64'hFFFFF7D5FFFFF7D5;
defparam \av_waitrequest~0 .shared_arith = "off";

cyclonev_lcell_comb \read_accepted~0 (
	.dataa(!clr_break_line),
	.datab(!d_read),
	.datac(!read_accepted1),
	.datad(!WideOr1),
	.datae(!WideOr0),
	.dataf(!WideOr01),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_accepted~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_accepted~0 .extended_lut = "off";
defparam \read_accepted~0 .lut_mask = 64'hFFFFFFFFFFFF7FFF;
defparam \read_accepted~0 .shared_arith = "off";

endmodule

module first_nios2_system_altera_merlin_slave_agent (
	mem_used_1,
	always1,
	m0_write)/* synthesis synthesis_greybox=1 */;
input 	mem_used_1;
input 	always1;
output 	m0_write;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \m0_write~0 (
	.dataa(!mem_used_1),
	.datab(!always1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(m0_write),
	.sumout(),
	.cout(),
	.shareout());
defparam \m0_write~0 .extended_lut = "off";
defparam \m0_write~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \m0_write~0 .shared_arith = "off";

endmodule

module first_nios2_system_altera_merlin_slave_agent_1 (
	always1,
	mem_used_1,
	m0_write)/* synthesis synthesis_greybox=1 */;
input 	always1;
input 	mem_used_1;
output 	m0_write;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \m0_write~0 (
	.dataa(!always1),
	.datab(!mem_used_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(m0_write),
	.sumout(),
	.cout(),
	.shareout());
defparam \m0_write~0 .extended_lut = "off";
defparam \m0_write~0 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \m0_write~0 .shared_arith = "off";

endmodule

module first_nios2_system_altera_merlin_slave_agent_2 (
	Equal6,
	always1,
	mem_used_1,
	m0_write)/* synthesis synthesis_greybox=1 */;
input 	Equal6;
input 	always1;
input 	mem_used_1;
output 	m0_write;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \m0_write~0 (
	.dataa(!Equal6),
	.datab(!always1),
	.datac(!mem_used_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(m0_write),
	.sumout(),
	.cout(),
	.shareout());
defparam \m0_write~0 .extended_lut = "off";
defparam \m0_write~0 .lut_mask = 64'hF7F7F7F7F7F7F7F7;
defparam \m0_write~0 .shared_arith = "off";

endmodule

module first_nios2_system_altera_merlin_slave_agent_3 (
	always1,
	mem_used_1,
	always11,
	m0_write)/* synthesis synthesis_greybox=1 */;
input 	always1;
input 	mem_used_1;
input 	always11;
output 	m0_write;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \m0_write~0 (
	.dataa(!always1),
	.datab(!mem_used_1),
	.datac(!always11),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(m0_write),
	.sumout(),
	.cout(),
	.shareout());
defparam \m0_write~0 .extended_lut = "off";
defparam \m0_write~0 .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \m0_write~0 .shared_arith = "off";

endmodule

module first_nios2_system_altera_merlin_slave_agent_6 (
	A_mem_baddr_5,
	A_mem_baddr_8,
	Equal1,
	Equal2,
	mem_used_1,
	Equal14,
	m0_write)/* synthesis synthesis_greybox=1 */;
input 	A_mem_baddr_5;
input 	A_mem_baddr_8;
input 	Equal1;
input 	Equal2;
input 	mem_used_1;
input 	Equal14;
output 	m0_write;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \m0_write~0 (
	.dataa(!A_mem_baddr_5),
	.datab(!A_mem_baddr_8),
	.datac(!Equal1),
	.datad(!Equal2),
	.datae(!mem_used_1),
	.dataf(!Equal14),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(m0_write),
	.sumout(),
	.cout(),
	.shareout());
defparam \m0_write~0 .extended_lut = "off";
defparam \m0_write~0 .lut_mask = 64'hFFFFEFFFFFFFFFFF;
defparam \m0_write~0 .shared_arith = "off";

endmodule

module first_nios2_system_altera_merlin_slave_agent_7 (
	mem_used_1,
	Equal6,
	m0_write)/* synthesis synthesis_greybox=1 */;
input 	mem_used_1;
input 	Equal6;
output 	m0_write;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \m0_write~0 (
	.dataa(!mem_used_1),
	.datab(!Equal6),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(m0_write),
	.sumout(),
	.cout(),
	.shareout());
defparam \m0_write~0 .extended_lut = "off";
defparam \m0_write~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \m0_write~0 .shared_arith = "off";

endmodule

module first_nios2_system_altera_merlin_slave_agent_8 (
	A_mem_baddr_7,
	mem_used_1,
	always1,
	m0_write)/* synthesis synthesis_greybox=1 */;
input 	A_mem_baddr_7;
input 	mem_used_1;
input 	always1;
output 	m0_write;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \m0_write~0 (
	.dataa(!A_mem_baddr_7),
	.datab(!mem_used_1),
	.datac(!always1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(m0_write),
	.sumout(),
	.cout(),
	.shareout());
defparam \m0_write~0 .extended_lut = "off";
defparam \m0_write~0 .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \m0_write~0 .shared_arith = "off";

endmodule

module first_nios2_system_altera_merlin_slave_agent_10 (
	mem_used_1,
	Equal16,
	m0_write)/* synthesis synthesis_greybox=1 */;
input 	mem_used_1;
input 	Equal16;
output 	m0_write;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \m0_write~0 (
	.dataa(!mem_used_1),
	.datab(!Equal16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(m0_write),
	.sumout(),
	.cout(),
	.shareout());
defparam \m0_write~0 .extended_lut = "off";
defparam \m0_write~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \m0_write~0 .shared_arith = "off";

endmodule

module first_nios2_system_altera_merlin_slave_agent_12 (
	mem_used_1,
	always1,
	m0_write)/* synthesis synthesis_greybox=1 */;
input 	mem_used_1;
input 	always1;
output 	m0_write;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \m0_write~0 (
	.dataa(!mem_used_1),
	.datab(!always1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(m0_write),
	.sumout(),
	.cout(),
	.shareout());
defparam \m0_write~0 .extended_lut = "off";
defparam \m0_write~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \m0_write~0 .shared_arith = "off";

endmodule

module first_nios2_system_altera_merlin_slave_agent_13 (
	mem_used_1,
	always1,
	m0_write)/* synthesis synthesis_greybox=1 */;
input 	mem_used_1;
input 	always1;
output 	m0_write;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \m0_write~0 (
	.dataa(!mem_used_1),
	.datab(!always1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(m0_write),
	.sumout(),
	.cout(),
	.shareout());
defparam \m0_write~0 .extended_lut = "off";
defparam \m0_write~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \m0_write~0 .shared_arith = "off";

endmodule

module first_nios2_system_altera_merlin_slave_agent_14 (
	A_mem_baddr_4,
	A_mem_baddr_7,
	A_mem_baddr_6,
	Equal2,
	mem_used_1,
	m0_write)/* synthesis synthesis_greybox=1 */;
input 	A_mem_baddr_4;
input 	A_mem_baddr_7;
input 	A_mem_baddr_6;
input 	Equal2;
input 	mem_used_1;
output 	m0_write;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \m0_write~0 (
	.dataa(!A_mem_baddr_4),
	.datab(!A_mem_baddr_7),
	.datac(!A_mem_baddr_6),
	.datad(!Equal2),
	.datae(!mem_used_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(m0_write),
	.sumout(),
	.cout(),
	.shareout());
defparam \m0_write~0 .extended_lut = "off";
defparam \m0_write~0 .lut_mask = 64'hFFFFFBFFFFFFFBFF;
defparam \m0_write~0 .shared_arith = "off";

endmodule

module first_nios2_system_altera_merlin_slave_agent_15 (
	Equal2,
	mem_used_1,
	m0_write)/* synthesis synthesis_greybox=1 */;
input 	Equal2;
input 	mem_used_1;
output 	m0_write;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \m0_write~0 (
	.dataa(!Equal2),
	.datab(!mem_used_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(m0_write),
	.sumout(),
	.cout(),
	.shareout());
defparam \m0_write~0 .extended_lut = "off";
defparam \m0_write~0 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \m0_write~0 .shared_arith = "off";

endmodule

module first_nios2_system_altera_merlin_slave_agent_17 (
	always1,
	mem_used_1,
	m0_write)/* synthesis synthesis_greybox=1 */;
input 	always1;
input 	mem_used_1;
output 	m0_write;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \m0_write~0 (
	.dataa(!always1),
	.datab(!mem_used_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(m0_write),
	.sumout(),
	.cout(),
	.shareout());
defparam \m0_write~0 .extended_lut = "off";
defparam \m0_write~0 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \m0_write~0 .shared_arith = "off";

endmodule

module first_nios2_system_altera_merlin_slave_agent_18 (
	clr_break_line,
	d_write,
	m0_write,
	always1,
	mem_used_1,
	m0_write1)/* synthesis synthesis_greybox=1 */;
input 	clr_break_line;
input 	d_write;
output 	m0_write;
input 	always1;
input 	mem_used_1;
output 	m0_write1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \m0_write~0 (
	.dataa(!clr_break_line),
	.datab(!d_write),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(m0_write),
	.sumout(),
	.cout(),
	.shareout());
defparam \m0_write~0 .extended_lut = "off";
defparam \m0_write~0 .lut_mask = 64'h7777777777777777;
defparam \m0_write~0 .shared_arith = "off";

cyclonev_lcell_comb \m0_write~1 (
	.dataa(!always1),
	.datab(!mem_used_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(m0_write1),
	.sumout(),
	.cout(),
	.shareout());
defparam \m0_write~1 .extended_lut = "off";
defparam \m0_write~1 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \m0_write~1 .shared_arith = "off";

endmodule

module first_nios2_system_altera_merlin_slave_translator (
	av_readdata,
	d_write,
	reset,
	cp_valid,
	read_latency_shift_reg_0,
	wait_latency_counter_1,
	wait_latency_counter_0,
	sink_ready,
	m0_write,
	av_readdata_pre_0,
	av_readdata_pre_1,
	av_readdata_pre_2,
	av_readdata_pre_3,
	av_readdata_pre_4,
	av_readdata_pre_5,
	av_readdata_pre_6,
	clk)/* synthesis synthesis_greybox=1 */;
input 	[31:0] av_readdata;
input 	d_write;
input 	reset;
input 	cp_valid;
output 	read_latency_shift_reg_0;
output 	wait_latency_counter_1;
output 	wait_latency_counter_0;
input 	sink_ready;
input 	m0_write;
output 	av_readdata_pre_0;
output 	av_readdata_pre_1;
output 	av_readdata_pre_2;
output 	av_readdata_pre_3;
output 	av_readdata_pre_4;
output 	av_readdata_pre_5;
output 	av_readdata_pre_6;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wait_latency_counter~0_combout ;
wire \wait_latency_counter~1_combout ;


dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(sink_ready),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

dffeas \wait_latency_counter[1] (
	.clk(clk),
	.d(\wait_latency_counter~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_1),
	.prn(vcc));
defparam \wait_latency_counter[1] .is_wysiwyg = "true";
defparam \wait_latency_counter[1] .power_up = "low";

dffeas \wait_latency_counter[0] (
	.clk(clk),
	.d(\wait_latency_counter~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_0),
	.prn(vcc));
defparam \wait_latency_counter[0] .is_wysiwyg = "true";
defparam \wait_latency_counter[0] .power_up = "low";

dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

dffeas \av_readdata_pre[1] (
	.clk(clk),
	.d(av_readdata[1]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_1),
	.prn(vcc));
defparam \av_readdata_pre[1] .is_wysiwyg = "true";
defparam \av_readdata_pre[1] .power_up = "low";

dffeas \av_readdata_pre[2] (
	.clk(clk),
	.d(av_readdata[2]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_2),
	.prn(vcc));
defparam \av_readdata_pre[2] .is_wysiwyg = "true";
defparam \av_readdata_pre[2] .power_up = "low";

dffeas \av_readdata_pre[3] (
	.clk(clk),
	.d(av_readdata[3]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_3),
	.prn(vcc));
defparam \av_readdata_pre[3] .is_wysiwyg = "true";
defparam \av_readdata_pre[3] .power_up = "low";

dffeas \av_readdata_pre[4] (
	.clk(clk),
	.d(av_readdata[4]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_4),
	.prn(vcc));
defparam \av_readdata_pre[4] .is_wysiwyg = "true";
defparam \av_readdata_pre[4] .power_up = "low";

dffeas \av_readdata_pre[5] (
	.clk(clk),
	.d(av_readdata[5]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_5),
	.prn(vcc));
defparam \av_readdata_pre[5] .is_wysiwyg = "true";
defparam \av_readdata_pre[5] .power_up = "low";

dffeas \av_readdata_pre[6] (
	.clk(clk),
	.d(av_readdata[6]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_6),
	.prn(vcc));
defparam \av_readdata_pre[6] .is_wysiwyg = "true";
defparam \av_readdata_pre[6] .power_up = "low";

cyclonev_lcell_comb \wait_latency_counter~0 (
	.dataa(!d_write),
	.datab(!cp_valid),
	.datac(!wait_latency_counter_1),
	.datad(!wait_latency_counter_0),
	.datae(!m0_write),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~0 .extended_lut = "off";
defparam \wait_latency_counter~0 .lut_mask = 64'h7FF7FFFF7FF7FFFF;
defparam \wait_latency_counter~0 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter~1 (
	.dataa(!d_write),
	.datab(!cp_valid),
	.datac(!wait_latency_counter_1),
	.datad(!wait_latency_counter_0),
	.datae(!m0_write),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~1 .extended_lut = "off";
defparam \wait_latency_counter~1 .lut_mask = 64'hFFBFFFFFFFBFFFFF;
defparam \wait_latency_counter~1 .shared_arith = "off";

endmodule

module first_nios2_system_altera_merlin_slave_translator_1 (
	av_readdata,
	d_write,
	reset,
	cp_valid,
	read_latency_shift_reg_0,
	wait_latency_counter_1,
	wait_latency_counter_0,
	sink_ready,
	m0_write,
	av_readdata_pre_0,
	av_readdata_pre_1,
	av_readdata_pre_2,
	av_readdata_pre_3,
	av_readdata_pre_4,
	av_readdata_pre_5,
	av_readdata_pre_6,
	clk)/* synthesis synthesis_greybox=1 */;
input 	[31:0] av_readdata;
input 	d_write;
input 	reset;
input 	cp_valid;
output 	read_latency_shift_reg_0;
output 	wait_latency_counter_1;
output 	wait_latency_counter_0;
input 	sink_ready;
input 	m0_write;
output 	av_readdata_pre_0;
output 	av_readdata_pre_1;
output 	av_readdata_pre_2;
output 	av_readdata_pre_3;
output 	av_readdata_pre_4;
output 	av_readdata_pre_5;
output 	av_readdata_pre_6;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wait_latency_counter~0_combout ;
wire \wait_latency_counter~1_combout ;


dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(sink_ready),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

dffeas \wait_latency_counter[1] (
	.clk(clk),
	.d(\wait_latency_counter~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_1),
	.prn(vcc));
defparam \wait_latency_counter[1] .is_wysiwyg = "true";
defparam \wait_latency_counter[1] .power_up = "low";

dffeas \wait_latency_counter[0] (
	.clk(clk),
	.d(\wait_latency_counter~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_0),
	.prn(vcc));
defparam \wait_latency_counter[0] .is_wysiwyg = "true";
defparam \wait_latency_counter[0] .power_up = "low";

dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

dffeas \av_readdata_pre[1] (
	.clk(clk),
	.d(av_readdata[1]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_1),
	.prn(vcc));
defparam \av_readdata_pre[1] .is_wysiwyg = "true";
defparam \av_readdata_pre[1] .power_up = "low";

dffeas \av_readdata_pre[2] (
	.clk(clk),
	.d(av_readdata[2]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_2),
	.prn(vcc));
defparam \av_readdata_pre[2] .is_wysiwyg = "true";
defparam \av_readdata_pre[2] .power_up = "low";

dffeas \av_readdata_pre[3] (
	.clk(clk),
	.d(av_readdata[3]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_3),
	.prn(vcc));
defparam \av_readdata_pre[3] .is_wysiwyg = "true";
defparam \av_readdata_pre[3] .power_up = "low";

dffeas \av_readdata_pre[4] (
	.clk(clk),
	.d(av_readdata[4]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_4),
	.prn(vcc));
defparam \av_readdata_pre[4] .is_wysiwyg = "true";
defparam \av_readdata_pre[4] .power_up = "low";

dffeas \av_readdata_pre[5] (
	.clk(clk),
	.d(av_readdata[5]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_5),
	.prn(vcc));
defparam \av_readdata_pre[5] .is_wysiwyg = "true";
defparam \av_readdata_pre[5] .power_up = "low";

dffeas \av_readdata_pre[6] (
	.clk(clk),
	.d(av_readdata[6]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_6),
	.prn(vcc));
defparam \av_readdata_pre[6] .is_wysiwyg = "true";
defparam \av_readdata_pre[6] .power_up = "low";

cyclonev_lcell_comb \wait_latency_counter~0 (
	.dataa(!d_write),
	.datab(!cp_valid),
	.datac(!wait_latency_counter_1),
	.datad(!wait_latency_counter_0),
	.datae(!m0_write),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~0 .extended_lut = "off";
defparam \wait_latency_counter~0 .lut_mask = 64'h7FF7FFFF7FF7FFFF;
defparam \wait_latency_counter~0 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter~1 (
	.dataa(!d_write),
	.datab(!cp_valid),
	.datac(!wait_latency_counter_1),
	.datad(!wait_latency_counter_0),
	.datae(!m0_write),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~1 .extended_lut = "off";
defparam \wait_latency_counter~1 .lut_mask = 64'hFFBFFFFFFFBFFFFF;
defparam \wait_latency_counter~1 .shared_arith = "off";

endmodule

module first_nios2_system_altera_merlin_slave_translator_2 (
	av_readdata,
	d_write,
	reset,
	Equal6,
	m0_write,
	cp_valid,
	read_latency_shift_reg_0,
	always1,
	mem_used_1,
	av_waitrequest_generated,
	sink_ready,
	m0_write1,
	av_readdata_pre_0,
	av_readdata_pre_1,
	av_readdata_pre_2,
	av_readdata_pre_3,
	av_readdata_pre_4,
	av_readdata_pre_5,
	clk)/* synthesis synthesis_greybox=1 */;
input 	[31:0] av_readdata;
input 	d_write;
input 	reset;
input 	Equal6;
input 	m0_write;
input 	cp_valid;
output 	read_latency_shift_reg_0;
input 	always1;
input 	mem_used_1;
output 	av_waitrequest_generated;
input 	sink_ready;
input 	m0_write1;
output 	av_readdata_pre_0;
output 	av_readdata_pre_1;
output 	av_readdata_pre_2;
output 	av_readdata_pre_3;
output 	av_readdata_pre_4;
output 	av_readdata_pre_5;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wait_latency_counter~1_combout ;
wire \wait_latency_counter[0]~q ;
wire \wait_latency_counter~0_combout ;
wire \wait_latency_counter[1]~q ;


dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(sink_ready),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

cyclonev_lcell_comb \av_waitrequest_generated~0 (
	.dataa(!Equal6),
	.datab(!m0_write),
	.datac(!always1),
	.datad(!mem_used_1),
	.datae(!\wait_latency_counter[1]~q ),
	.dataf(!\wait_latency_counter[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(av_waitrequest_generated),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_waitrequest_generated~0 .extended_lut = "off";
defparam \av_waitrequest_generated~0 .lut_mask = 64'hFFFF9669FFFF6996;
defparam \av_waitrequest_generated~0 .shared_arith = "off";

dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

dffeas \av_readdata_pre[1] (
	.clk(clk),
	.d(av_readdata[1]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_1),
	.prn(vcc));
defparam \av_readdata_pre[1] .is_wysiwyg = "true";
defparam \av_readdata_pre[1] .power_up = "low";

dffeas \av_readdata_pre[2] (
	.clk(clk),
	.d(av_readdata[2]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_2),
	.prn(vcc));
defparam \av_readdata_pre[2] .is_wysiwyg = "true";
defparam \av_readdata_pre[2] .power_up = "low";

dffeas \av_readdata_pre[3] (
	.clk(clk),
	.d(av_readdata[3]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_3),
	.prn(vcc));
defparam \av_readdata_pre[3] .is_wysiwyg = "true";
defparam \av_readdata_pre[3] .power_up = "low";

dffeas \av_readdata_pre[4] (
	.clk(clk),
	.d(av_readdata[4]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_4),
	.prn(vcc));
defparam \av_readdata_pre[4] .is_wysiwyg = "true";
defparam \av_readdata_pre[4] .power_up = "low";

dffeas \av_readdata_pre[5] (
	.clk(clk),
	.d(av_readdata[5]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_5),
	.prn(vcc));
defparam \av_readdata_pre[5] .is_wysiwyg = "true";
defparam \av_readdata_pre[5] .power_up = "low";

cyclonev_lcell_comb \wait_latency_counter~1 (
	.dataa(!cp_valid),
	.datab(!\wait_latency_counter[0]~q ),
	.datac(!m0_write1),
	.datad(!av_waitrequest_generated),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~1 .extended_lut = "off";
defparam \wait_latency_counter~1 .lut_mask = 64'hFFDFFFDFFFDFFFDF;
defparam \wait_latency_counter~1 .shared_arith = "off";

dffeas \wait_latency_counter[0] (
	.clk(clk),
	.d(\wait_latency_counter~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wait_latency_counter[0]~q ),
	.prn(vcc));
defparam \wait_latency_counter[0] .is_wysiwyg = "true";
defparam \wait_latency_counter[0] .power_up = "low";

cyclonev_lcell_comb \wait_latency_counter~0 (
	.dataa(!d_write),
	.datab(!cp_valid),
	.datac(!\wait_latency_counter[1]~q ),
	.datad(!\wait_latency_counter[0]~q ),
	.datae(!m0_write1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~0 .extended_lut = "off";
defparam \wait_latency_counter~0 .lut_mask = 64'h7FF7FFFF7FF7FFFF;
defparam \wait_latency_counter~0 .shared_arith = "off";

dffeas \wait_latency_counter[1] (
	.clk(clk),
	.d(\wait_latency_counter~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wait_latency_counter[1]~q ),
	.prn(vcc));
defparam \wait_latency_counter[1] .is_wysiwyg = "true";
defparam \wait_latency_counter[1] .power_up = "low";

endmodule

module first_nios2_system_altera_merlin_slave_translator_3 (
	av_readdata,
	d_write,
	reset,
	m0_write,
	cp_valid,
	read_latency_shift_reg_0,
	always1,
	mem_used_1,
	always11,
	av_waitrequest_generated,
	sink_ready,
	m0_write1,
	av_readdata_pre_0,
	av_readdata_pre_1,
	av_readdata_pre_2,
	av_readdata_pre_3,
	av_readdata_pre_4,
	av_readdata_pre_5,
	clk)/* synthesis synthesis_greybox=1 */;
input 	[31:0] av_readdata;
input 	d_write;
input 	reset;
input 	m0_write;
input 	cp_valid;
output 	read_latency_shift_reg_0;
input 	always1;
input 	mem_used_1;
input 	always11;
output 	av_waitrequest_generated;
input 	sink_ready;
input 	m0_write1;
output 	av_readdata_pre_0;
output 	av_readdata_pre_1;
output 	av_readdata_pre_2;
output 	av_readdata_pre_3;
output 	av_readdata_pre_4;
output 	av_readdata_pre_5;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wait_latency_counter~1_combout ;
wire \wait_latency_counter[0]~q ;
wire \wait_latency_counter~0_combout ;
wire \wait_latency_counter[1]~q ;


dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(sink_ready),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

cyclonev_lcell_comb \av_waitrequest_generated~0 (
	.dataa(!m0_write),
	.datab(!always1),
	.datac(!mem_used_1),
	.datad(!\wait_latency_counter[1]~q ),
	.datae(!\wait_latency_counter[0]~q ),
	.dataf(!always11),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(av_waitrequest_generated),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_waitrequest_generated~0 .extended_lut = "off";
defparam \av_waitrequest_generated~0 .lut_mask = 64'hFF96FF69FF69FF96;
defparam \av_waitrequest_generated~0 .shared_arith = "off";

dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

dffeas \av_readdata_pre[1] (
	.clk(clk),
	.d(av_readdata[1]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_1),
	.prn(vcc));
defparam \av_readdata_pre[1] .is_wysiwyg = "true";
defparam \av_readdata_pre[1] .power_up = "low";

dffeas \av_readdata_pre[2] (
	.clk(clk),
	.d(av_readdata[2]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_2),
	.prn(vcc));
defparam \av_readdata_pre[2] .is_wysiwyg = "true";
defparam \av_readdata_pre[2] .power_up = "low";

dffeas \av_readdata_pre[3] (
	.clk(clk),
	.d(av_readdata[3]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_3),
	.prn(vcc));
defparam \av_readdata_pre[3] .is_wysiwyg = "true";
defparam \av_readdata_pre[3] .power_up = "low";

dffeas \av_readdata_pre[4] (
	.clk(clk),
	.d(av_readdata[4]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_4),
	.prn(vcc));
defparam \av_readdata_pre[4] .is_wysiwyg = "true";
defparam \av_readdata_pre[4] .power_up = "low";

dffeas \av_readdata_pre[5] (
	.clk(clk),
	.d(av_readdata[5]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_5),
	.prn(vcc));
defparam \av_readdata_pre[5] .is_wysiwyg = "true";
defparam \av_readdata_pre[5] .power_up = "low";

cyclonev_lcell_comb \wait_latency_counter~1 (
	.dataa(!cp_valid),
	.datab(!\wait_latency_counter[0]~q ),
	.datac(!m0_write1),
	.datad(!av_waitrequest_generated),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~1 .extended_lut = "off";
defparam \wait_latency_counter~1 .lut_mask = 64'hFFDFFFDFFFDFFFDF;
defparam \wait_latency_counter~1 .shared_arith = "off";

dffeas \wait_latency_counter[0] (
	.clk(clk),
	.d(\wait_latency_counter~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wait_latency_counter[0]~q ),
	.prn(vcc));
defparam \wait_latency_counter[0] .is_wysiwyg = "true";
defparam \wait_latency_counter[0] .power_up = "low";

cyclonev_lcell_comb \wait_latency_counter~0 (
	.dataa(!d_write),
	.datab(!cp_valid),
	.datac(!\wait_latency_counter[1]~q ),
	.datad(!\wait_latency_counter[0]~q ),
	.datae(!m0_write1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~0 .extended_lut = "off";
defparam \wait_latency_counter~0 .lut_mask = 64'h7FF7FFFF7FF7FFFF;
defparam \wait_latency_counter~0 .shared_arith = "off";

dffeas \wait_latency_counter[1] (
	.clk(clk),
	.d(\wait_latency_counter~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wait_latency_counter[1]~q ),
	.prn(vcc));
defparam \wait_latency_counter[1] .is_wysiwyg = "true";
defparam \wait_latency_counter[1] .power_up = "low";

endmodule

module first_nios2_system_altera_merlin_slave_translator_4 (
	av_readdata,
	clr_break_line,
	reset,
	read_latency_shift_reg_0,
	write,
	WideOr1,
	mem,
	av_readdata_pre_0,
	av_readdata_pre_1,
	av_readdata_pre_2,
	av_readdata_pre_3,
	av_readdata_pre_4,
	av_readdata_pre_5,
	av_readdata_pre_6,
	av_readdata_pre_7,
	av_readdata_pre_22,
	av_readdata_pre_23,
	av_readdata_pre_24,
	av_readdata_pre_25,
	av_readdata_pre_31,
	av_readdata_pre_21,
	av_readdata_pre_11,
	av_readdata_pre_28,
	av_readdata_pre_10,
	av_readdata_pre_27,
	av_readdata_pre_8,
	av_readdata_pre_9,
	av_readdata_pre_26,
	av_readdata_pre_20,
	av_readdata_pre_19,
	av_readdata_pre_17,
	av_readdata_pre_30,
	av_readdata_pre_18,
	av_readdata_pre_16,
	av_readdata_pre_15,
	av_readdata_pre_12,
	av_readdata_pre_13,
	av_readdata_pre_14,
	av_readdata_pre_29,
	clk)/* synthesis synthesis_greybox=1 */;
input 	[31:0] av_readdata;
input 	clr_break_line;
input 	reset;
output 	read_latency_shift_reg_0;
input 	write;
input 	WideOr1;
input 	mem;
output 	av_readdata_pre_0;
output 	av_readdata_pre_1;
output 	av_readdata_pre_2;
output 	av_readdata_pre_3;
output 	av_readdata_pre_4;
output 	av_readdata_pre_5;
output 	av_readdata_pre_6;
output 	av_readdata_pre_7;
output 	av_readdata_pre_22;
output 	av_readdata_pre_23;
output 	av_readdata_pre_24;
output 	av_readdata_pre_25;
output 	av_readdata_pre_31;
output 	av_readdata_pre_21;
output 	av_readdata_pre_11;
output 	av_readdata_pre_28;
output 	av_readdata_pre_10;
output 	av_readdata_pre_27;
output 	av_readdata_pre_8;
output 	av_readdata_pre_9;
output 	av_readdata_pre_26;
output 	av_readdata_pre_20;
output 	av_readdata_pre_19;
output 	av_readdata_pre_17;
output 	av_readdata_pre_30;
output 	av_readdata_pre_18;
output 	av_readdata_pre_16;
output 	av_readdata_pre_15;
output 	av_readdata_pre_12;
output 	av_readdata_pre_13;
output 	av_readdata_pre_14;
output 	av_readdata_pre_29;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read_latency_shift_reg~0_combout ;


dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(\read_latency_shift_reg~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

dffeas \av_readdata_pre[1] (
	.clk(clk),
	.d(av_readdata[1]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_1),
	.prn(vcc));
defparam \av_readdata_pre[1] .is_wysiwyg = "true";
defparam \av_readdata_pre[1] .power_up = "low";

dffeas \av_readdata_pre[2] (
	.clk(clk),
	.d(av_readdata[2]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_2),
	.prn(vcc));
defparam \av_readdata_pre[2] .is_wysiwyg = "true";
defparam \av_readdata_pre[2] .power_up = "low";

dffeas \av_readdata_pre[3] (
	.clk(clk),
	.d(av_readdata[3]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_3),
	.prn(vcc));
defparam \av_readdata_pre[3] .is_wysiwyg = "true";
defparam \av_readdata_pre[3] .power_up = "low";

dffeas \av_readdata_pre[4] (
	.clk(clk),
	.d(av_readdata[4]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_4),
	.prn(vcc));
defparam \av_readdata_pre[4] .is_wysiwyg = "true";
defparam \av_readdata_pre[4] .power_up = "low";

dffeas \av_readdata_pre[5] (
	.clk(clk),
	.d(av_readdata[5]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_5),
	.prn(vcc));
defparam \av_readdata_pre[5] .is_wysiwyg = "true";
defparam \av_readdata_pre[5] .power_up = "low";

dffeas \av_readdata_pre[6] (
	.clk(clk),
	.d(av_readdata[6]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_6),
	.prn(vcc));
defparam \av_readdata_pre[6] .is_wysiwyg = "true";
defparam \av_readdata_pre[6] .power_up = "low";

dffeas \av_readdata_pre[7] (
	.clk(clk),
	.d(av_readdata[7]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_7),
	.prn(vcc));
defparam \av_readdata_pre[7] .is_wysiwyg = "true";
defparam \av_readdata_pre[7] .power_up = "low";

dffeas \av_readdata_pre[22] (
	.clk(clk),
	.d(av_readdata[22]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_22),
	.prn(vcc));
defparam \av_readdata_pre[22] .is_wysiwyg = "true";
defparam \av_readdata_pre[22] .power_up = "low";

dffeas \av_readdata_pre[23] (
	.clk(clk),
	.d(av_readdata[23]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_23),
	.prn(vcc));
defparam \av_readdata_pre[23] .is_wysiwyg = "true";
defparam \av_readdata_pre[23] .power_up = "low";

dffeas \av_readdata_pre[24] (
	.clk(clk),
	.d(av_readdata[24]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_24),
	.prn(vcc));
defparam \av_readdata_pre[24] .is_wysiwyg = "true";
defparam \av_readdata_pre[24] .power_up = "low";

dffeas \av_readdata_pre[25] (
	.clk(clk),
	.d(av_readdata[25]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_25),
	.prn(vcc));
defparam \av_readdata_pre[25] .is_wysiwyg = "true";
defparam \av_readdata_pre[25] .power_up = "low";

dffeas \av_readdata_pre[31] (
	.clk(clk),
	.d(av_readdata[31]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_31),
	.prn(vcc));
defparam \av_readdata_pre[31] .is_wysiwyg = "true";
defparam \av_readdata_pre[31] .power_up = "low";

dffeas \av_readdata_pre[21] (
	.clk(clk),
	.d(av_readdata[21]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_21),
	.prn(vcc));
defparam \av_readdata_pre[21] .is_wysiwyg = "true";
defparam \av_readdata_pre[21] .power_up = "low";

dffeas \av_readdata_pre[11] (
	.clk(clk),
	.d(av_readdata[11]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_11),
	.prn(vcc));
defparam \av_readdata_pre[11] .is_wysiwyg = "true";
defparam \av_readdata_pre[11] .power_up = "low";

dffeas \av_readdata_pre[28] (
	.clk(clk),
	.d(av_readdata[28]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_28),
	.prn(vcc));
defparam \av_readdata_pre[28] .is_wysiwyg = "true";
defparam \av_readdata_pre[28] .power_up = "low";

dffeas \av_readdata_pre[10] (
	.clk(clk),
	.d(av_readdata[10]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_10),
	.prn(vcc));
defparam \av_readdata_pre[10] .is_wysiwyg = "true";
defparam \av_readdata_pre[10] .power_up = "low";

dffeas \av_readdata_pre[27] (
	.clk(clk),
	.d(av_readdata[27]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_27),
	.prn(vcc));
defparam \av_readdata_pre[27] .is_wysiwyg = "true";
defparam \av_readdata_pre[27] .power_up = "low";

dffeas \av_readdata_pre[8] (
	.clk(clk),
	.d(av_readdata[8]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_8),
	.prn(vcc));
defparam \av_readdata_pre[8] .is_wysiwyg = "true";
defparam \av_readdata_pre[8] .power_up = "low";

dffeas \av_readdata_pre[9] (
	.clk(clk),
	.d(av_readdata[9]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_9),
	.prn(vcc));
defparam \av_readdata_pre[9] .is_wysiwyg = "true";
defparam \av_readdata_pre[9] .power_up = "low";

dffeas \av_readdata_pre[26] (
	.clk(clk),
	.d(av_readdata[26]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_26),
	.prn(vcc));
defparam \av_readdata_pre[26] .is_wysiwyg = "true";
defparam \av_readdata_pre[26] .power_up = "low";

dffeas \av_readdata_pre[20] (
	.clk(clk),
	.d(av_readdata[20]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_20),
	.prn(vcc));
defparam \av_readdata_pre[20] .is_wysiwyg = "true";
defparam \av_readdata_pre[20] .power_up = "low";

dffeas \av_readdata_pre[19] (
	.clk(clk),
	.d(av_readdata[19]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_19),
	.prn(vcc));
defparam \av_readdata_pre[19] .is_wysiwyg = "true";
defparam \av_readdata_pre[19] .power_up = "low";

dffeas \av_readdata_pre[17] (
	.clk(clk),
	.d(av_readdata[17]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_17),
	.prn(vcc));
defparam \av_readdata_pre[17] .is_wysiwyg = "true";
defparam \av_readdata_pre[17] .power_up = "low";

dffeas \av_readdata_pre[30] (
	.clk(clk),
	.d(av_readdata[30]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_30),
	.prn(vcc));
defparam \av_readdata_pre[30] .is_wysiwyg = "true";
defparam \av_readdata_pre[30] .power_up = "low";

dffeas \av_readdata_pre[18] (
	.clk(clk),
	.d(av_readdata[18]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_18),
	.prn(vcc));
defparam \av_readdata_pre[18] .is_wysiwyg = "true";
defparam \av_readdata_pre[18] .power_up = "low";

dffeas \av_readdata_pre[16] (
	.clk(clk),
	.d(av_readdata[16]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_16),
	.prn(vcc));
defparam \av_readdata_pre[16] .is_wysiwyg = "true";
defparam \av_readdata_pre[16] .power_up = "low";

dffeas \av_readdata_pre[15] (
	.clk(clk),
	.d(av_readdata[15]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_15),
	.prn(vcc));
defparam \av_readdata_pre[15] .is_wysiwyg = "true";
defparam \av_readdata_pre[15] .power_up = "low";

dffeas \av_readdata_pre[12] (
	.clk(clk),
	.d(av_readdata[12]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_12),
	.prn(vcc));
defparam \av_readdata_pre[12] .is_wysiwyg = "true";
defparam \av_readdata_pre[12] .power_up = "low";

dffeas \av_readdata_pre[13] (
	.clk(clk),
	.d(av_readdata[13]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_13),
	.prn(vcc));
defparam \av_readdata_pre[13] .is_wysiwyg = "true";
defparam \av_readdata_pre[13] .power_up = "low";

dffeas \av_readdata_pre[14] (
	.clk(clk),
	.d(av_readdata[14]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_14),
	.prn(vcc));
defparam \av_readdata_pre[14] .is_wysiwyg = "true";
defparam \av_readdata_pre[14] .power_up = "low";

dffeas \av_readdata_pre[29] (
	.clk(clk),
	.d(av_readdata[29]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_29),
	.prn(vcc));
defparam \av_readdata_pre[29] .is_wysiwyg = "true";
defparam \av_readdata_pre[29] .power_up = "low";

cyclonev_lcell_comb \read_latency_shift_reg~0 (
	.dataa(!clr_break_line),
	.datab(!write),
	.datac(!WideOr1),
	.datad(!mem),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_latency_shift_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~0 .extended_lut = "off";
defparam \read_latency_shift_reg~0 .lut_mask = 64'hF7FFF7FFF7FFF7FF;
defparam \read_latency_shift_reg~0 .shared_arith = "off";

endmodule

module first_nios2_system_altera_merlin_slave_translator_5 (
	av_readdata_pre_0,
	av_readdata,
	always0,
	clr_break_line,
	wait_latency_counter_1,
	wait_latency_counter_0,
	d_write,
	Equal0,
	reset,
	read_latency_shift_reg_0,
	uav_read,
	read_latency_shift_reg,
	cp_valid,
	write,
	read_latency_shift_reg1,
	clk)/* synthesis synthesis_greybox=1 */;
output 	av_readdata_pre_0;
input 	[31:0] av_readdata;
input 	always0;
input 	clr_break_line;
output 	wait_latency_counter_1;
output 	wait_latency_counter_0;
input 	d_write;
input 	Equal0;
input 	reset;
output 	read_latency_shift_reg_0;
input 	uav_read;
output 	read_latency_shift_reg;
input 	cp_valid;
input 	write;
output 	read_latency_shift_reg1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wait_latency_counter~0_combout ;
wire \wait_latency_counter~1_combout ;


dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(Equal0),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

dffeas \wait_latency_counter[1] (
	.clk(clk),
	.d(\wait_latency_counter~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_1),
	.prn(vcc));
defparam \wait_latency_counter[1] .is_wysiwyg = "true";
defparam \wait_latency_counter[1] .power_up = "low";

dffeas \wait_latency_counter[0] (
	.clk(clk),
	.d(\wait_latency_counter~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_0),
	.prn(vcc));
defparam \wait_latency_counter[0] .is_wysiwyg = "true";
defparam \wait_latency_counter[0] .power_up = "low";

dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(read_latency_shift_reg1),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

cyclonev_lcell_comb \read_latency_shift_reg~0 (
	.dataa(!clr_break_line),
	.datab(!uav_read),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(read_latency_shift_reg),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~0 .extended_lut = "off";
defparam \read_latency_shift_reg~0 .lut_mask = 64'h7777777777777777;
defparam \read_latency_shift_reg~0 .shared_arith = "off";

cyclonev_lcell_comb \read_latency_shift_reg~1 (
	.dataa(!write),
	.datab(!read_latency_shift_reg),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(read_latency_shift_reg1),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~1 .extended_lut = "off";
defparam \read_latency_shift_reg~1 .lut_mask = 64'h7777777777777777;
defparam \read_latency_shift_reg~1 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter~0 (
	.dataa(!wait_latency_counter_1),
	.datab(!wait_latency_counter_0),
	.datac(!d_write),
	.datad(!always0),
	.datae(!cp_valid),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~0 .extended_lut = "off";
defparam \wait_latency_counter~0 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \wait_latency_counter~0 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter~1 (
	.dataa(!wait_latency_counter_1),
	.datab(!wait_latency_counter_0),
	.datac(!d_write),
	.datad(!always0),
	.datae(!cp_valid),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~1 .extended_lut = "off";
defparam \wait_latency_counter~1 .lut_mask = 64'hFDFFFFFFFDFFFFFF;
defparam \wait_latency_counter~1 .shared_arith = "off";

endmodule

module first_nios2_system_altera_merlin_slave_translator_6 (
	av_readdata_pre_0,
	av_readdata,
	clr_break_line,
	d_write,
	Equal0,
	reset,
	wait_latency_counter_1,
	m0_write,
	wait_latency_counter_0,
	uav_read,
	cp_valid,
	read_latency_shift_reg_0,
	clk)/* synthesis synthesis_greybox=1 */;
output 	av_readdata_pre_0;
input 	[31:0] av_readdata;
input 	clr_break_line;
input 	d_write;
input 	Equal0;
input 	reset;
output 	wait_latency_counter_1;
input 	m0_write;
output 	wait_latency_counter_0;
input 	uav_read;
input 	cp_valid;
output 	read_latency_shift_reg_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wait_latency_counter~0_combout ;
wire \wait_latency_counter~1_combout ;
wire \read_latency_shift_reg~0_combout ;


dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(Equal0),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

dffeas \wait_latency_counter[1] (
	.clk(clk),
	.d(\wait_latency_counter~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_1),
	.prn(vcc));
defparam \wait_latency_counter[1] .is_wysiwyg = "true";
defparam \wait_latency_counter[1] .power_up = "low";

dffeas \wait_latency_counter[0] (
	.clk(clk),
	.d(\wait_latency_counter~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_0),
	.prn(vcc));
defparam \wait_latency_counter[0] .is_wysiwyg = "true";
defparam \wait_latency_counter[0] .power_up = "low";

dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(\read_latency_shift_reg~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

cyclonev_lcell_comb \wait_latency_counter~0 (
	.dataa(!d_write),
	.datab(!wait_latency_counter_0),
	.datac(!wait_latency_counter_1),
	.datad(!m0_write),
	.datae(!cp_valid),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~0 .extended_lut = "off";
defparam \wait_latency_counter~0 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \wait_latency_counter~0 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter~1 (
	.dataa(!d_write),
	.datab(!wait_latency_counter_0),
	.datac(!wait_latency_counter_1),
	.datad(!m0_write),
	.datae(!cp_valid),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~1 .extended_lut = "off";
defparam \wait_latency_counter~1 .lut_mask = 64'hEFFFFFFFEFFFFFFF;
defparam \wait_latency_counter~1 .shared_arith = "off";

cyclonev_lcell_comb \read_latency_shift_reg~0 (
	.dataa(!clr_break_line),
	.datab(!d_write),
	.datac(!wait_latency_counter_0),
	.datad(!wait_latency_counter_1),
	.datae(!m0_write),
	.dataf(!uav_read),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_latency_shift_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~0 .extended_lut = "off";
defparam \read_latency_shift_reg~0 .lut_mask = 64'hFF7DFFFFFFFFFFFF;
defparam \read_latency_shift_reg~0 .shared_arith = "off";

endmodule

module first_nios2_system_altera_merlin_slave_translator_7 (
	av_readdata_pre_0,
	av_readdata_pre_1,
	av_readdata_pre_2,
	av_readdata_pre_3,
	av_readdata_pre_4,
	av_readdata_pre_5,
	av_readdata_pre_6,
	av_readdata,
	clr_break_line,
	d_write,
	Equal0,
	reset,
	wait_latency_counter_1,
	wait_latency_counter_0,
	m0_write,
	uav_read,
	cp_valid,
	read_latency_shift_reg_0,
	m0_write1,
	av_waitrequest_generated,
	clk)/* synthesis synthesis_greybox=1 */;
output 	av_readdata_pre_0;
output 	av_readdata_pre_1;
output 	av_readdata_pre_2;
output 	av_readdata_pre_3;
output 	av_readdata_pre_4;
output 	av_readdata_pre_5;
output 	av_readdata_pre_6;
input 	[31:0] av_readdata;
input 	clr_break_line;
input 	d_write;
input 	Equal0;
input 	reset;
output 	wait_latency_counter_1;
output 	wait_latency_counter_0;
input 	m0_write;
input 	uav_read;
input 	cp_valid;
output 	read_latency_shift_reg_0;
input 	m0_write1;
output 	av_waitrequest_generated;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wait_latency_counter~0_combout ;
wire \wait_latency_counter~1_combout ;
wire \read_latency_shift_reg~0_combout ;


dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(Equal0),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

dffeas \av_readdata_pre[1] (
	.clk(clk),
	.d(av_readdata[1]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(Equal0),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_1),
	.prn(vcc));
defparam \av_readdata_pre[1] .is_wysiwyg = "true";
defparam \av_readdata_pre[1] .power_up = "low";

dffeas \av_readdata_pre[2] (
	.clk(clk),
	.d(av_readdata[2]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(Equal0),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_2),
	.prn(vcc));
defparam \av_readdata_pre[2] .is_wysiwyg = "true";
defparam \av_readdata_pre[2] .power_up = "low";

dffeas \av_readdata_pre[3] (
	.clk(clk),
	.d(av_readdata[3]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(Equal0),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_3),
	.prn(vcc));
defparam \av_readdata_pre[3] .is_wysiwyg = "true";
defparam \av_readdata_pre[3] .power_up = "low";

dffeas \av_readdata_pre[4] (
	.clk(clk),
	.d(av_readdata[4]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(Equal0),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_4),
	.prn(vcc));
defparam \av_readdata_pre[4] .is_wysiwyg = "true";
defparam \av_readdata_pre[4] .power_up = "low";

dffeas \av_readdata_pre[5] (
	.clk(clk),
	.d(av_readdata[5]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(Equal0),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_5),
	.prn(vcc));
defparam \av_readdata_pre[5] .is_wysiwyg = "true";
defparam \av_readdata_pre[5] .power_up = "low";

dffeas \av_readdata_pre[6] (
	.clk(clk),
	.d(av_readdata[6]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(Equal0),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_6),
	.prn(vcc));
defparam \av_readdata_pre[6] .is_wysiwyg = "true";
defparam \av_readdata_pre[6] .power_up = "low";

dffeas \wait_latency_counter[1] (
	.clk(clk),
	.d(\wait_latency_counter~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_1),
	.prn(vcc));
defparam \wait_latency_counter[1] .is_wysiwyg = "true";
defparam \wait_latency_counter[1] .power_up = "low";

dffeas \wait_latency_counter[0] (
	.clk(clk),
	.d(\wait_latency_counter~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_0),
	.prn(vcc));
defparam \wait_latency_counter[0] .is_wysiwyg = "true";
defparam \wait_latency_counter[0] .power_up = "low";

dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(\read_latency_shift_reg~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

cyclonev_lcell_comb \av_waitrequest_generated~0 (
	.dataa(!wait_latency_counter_0),
	.datab(!wait_latency_counter_1),
	.datac(!m0_write1),
	.datad(!m0_write),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(av_waitrequest_generated),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_waitrequest_generated~0 .extended_lut = "off";
defparam \av_waitrequest_generated~0 .lut_mask = 64'hEDDEEDDEEDDEEDDE;
defparam \av_waitrequest_generated~0 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter~0 (
	.dataa(!d_write),
	.datab(!wait_latency_counter_0),
	.datac(!wait_latency_counter_1),
	.datad(!m0_write1),
	.datae(!cp_valid),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~0 .extended_lut = "off";
defparam \wait_latency_counter~0 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \wait_latency_counter~0 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter~1 (
	.dataa(!wait_latency_counter_0),
	.datab(!m0_write1),
	.datac(!cp_valid),
	.datad(!av_waitrequest_generated),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~1 .extended_lut = "off";
defparam \wait_latency_counter~1 .lut_mask = 64'hFFBFFFBFFFBFFFBF;
defparam \wait_latency_counter~1 .shared_arith = "off";

cyclonev_lcell_comb \read_latency_shift_reg~0 (
	.dataa(!clr_break_line),
	.datab(!d_write),
	.datac(!wait_latency_counter_0),
	.datad(!wait_latency_counter_1),
	.datae(!m0_write1),
	.dataf(!uav_read),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_latency_shift_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~0 .extended_lut = "off";
defparam \read_latency_shift_reg~0 .lut_mask = 64'hFF7DFFFFFFFFFFFF;
defparam \read_latency_shift_reg~0 .shared_arith = "off";

endmodule

module first_nios2_system_altera_merlin_slave_translator_8 (
	av_readdata_pre_0,
	av_readdata_pre_1,
	av_readdata_pre_2,
	av_readdata_pre_3,
	av_readdata_pre_4,
	av_readdata_pre_5,
	av_readdata_pre_6,
	av_readdata,
	A_mem_baddr_7,
	clr_break_line,
	d_write,
	Equal0,
	reset,
	wait_latency_counter_1,
	mem_used_1,
	always1,
	wait_latency_counter_0,
	m0_write,
	uav_read,
	cp_valid,
	read_latency_shift_reg_0,
	m0_write1,
	av_waitrequest_generated,
	clk)/* synthesis synthesis_greybox=1 */;
output 	av_readdata_pre_0;
output 	av_readdata_pre_1;
output 	av_readdata_pre_2;
output 	av_readdata_pre_3;
output 	av_readdata_pre_4;
output 	av_readdata_pre_5;
output 	av_readdata_pre_6;
input 	[31:0] av_readdata;
input 	A_mem_baddr_7;
input 	clr_break_line;
input 	d_write;
input 	Equal0;
input 	reset;
output 	wait_latency_counter_1;
input 	mem_used_1;
input 	always1;
output 	wait_latency_counter_0;
input 	m0_write;
input 	uav_read;
input 	cp_valid;
output 	read_latency_shift_reg_0;
input 	m0_write1;
output 	av_waitrequest_generated;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wait_latency_counter~0_combout ;
wire \wait_latency_counter~1_combout ;
wire \read_latency_shift_reg~0_combout ;


dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(Equal0),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

dffeas \av_readdata_pre[1] (
	.clk(clk),
	.d(av_readdata[1]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(Equal0),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_1),
	.prn(vcc));
defparam \av_readdata_pre[1] .is_wysiwyg = "true";
defparam \av_readdata_pre[1] .power_up = "low";

dffeas \av_readdata_pre[2] (
	.clk(clk),
	.d(av_readdata[2]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(Equal0),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_2),
	.prn(vcc));
defparam \av_readdata_pre[2] .is_wysiwyg = "true";
defparam \av_readdata_pre[2] .power_up = "low";

dffeas \av_readdata_pre[3] (
	.clk(clk),
	.d(av_readdata[3]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(Equal0),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_3),
	.prn(vcc));
defparam \av_readdata_pre[3] .is_wysiwyg = "true";
defparam \av_readdata_pre[3] .power_up = "low";

dffeas \av_readdata_pre[4] (
	.clk(clk),
	.d(av_readdata[4]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(Equal0),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_4),
	.prn(vcc));
defparam \av_readdata_pre[4] .is_wysiwyg = "true";
defparam \av_readdata_pre[4] .power_up = "low";

dffeas \av_readdata_pre[5] (
	.clk(clk),
	.d(av_readdata[5]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(Equal0),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_5),
	.prn(vcc));
defparam \av_readdata_pre[5] .is_wysiwyg = "true";
defparam \av_readdata_pre[5] .power_up = "low";

dffeas \av_readdata_pre[6] (
	.clk(clk),
	.d(av_readdata[6]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(Equal0),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_6),
	.prn(vcc));
defparam \av_readdata_pre[6] .is_wysiwyg = "true";
defparam \av_readdata_pre[6] .power_up = "low";

dffeas \wait_latency_counter[1] (
	.clk(clk),
	.d(\wait_latency_counter~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_1),
	.prn(vcc));
defparam \wait_latency_counter[1] .is_wysiwyg = "true";
defparam \wait_latency_counter[1] .power_up = "low";

dffeas \wait_latency_counter[0] (
	.clk(clk),
	.d(\wait_latency_counter~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_0),
	.prn(vcc));
defparam \wait_latency_counter[0] .is_wysiwyg = "true";
defparam \wait_latency_counter[0] .power_up = "low";

dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(\read_latency_shift_reg~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

cyclonev_lcell_comb \av_waitrequest_generated~0 (
	.dataa(!A_mem_baddr_7),
	.datab(!wait_latency_counter_0),
	.datac(!mem_used_1),
	.datad(!always1),
	.datae(!m0_write),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(av_waitrequest_generated),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_waitrequest_generated~0 .extended_lut = "off";
defparam \av_waitrequest_generated~0 .lut_mask = 64'h9669699696696996;
defparam \av_waitrequest_generated~0 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter~0 (
	.dataa(!d_write),
	.datab(!wait_latency_counter_0),
	.datac(!wait_latency_counter_1),
	.datad(!m0_write1),
	.datae(!cp_valid),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~0 .extended_lut = "off";
defparam \wait_latency_counter~0 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \wait_latency_counter~0 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter~1 (
	.dataa(!d_write),
	.datab(!wait_latency_counter_0),
	.datac(!wait_latency_counter_1),
	.datad(!m0_write1),
	.datae(!cp_valid),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~1 .extended_lut = "off";
defparam \wait_latency_counter~1 .lut_mask = 64'hEFFFFFFFEFFFFFFF;
defparam \wait_latency_counter~1 .shared_arith = "off";

cyclonev_lcell_comb \read_latency_shift_reg~0 (
	.dataa(!clr_break_line),
	.datab(!wait_latency_counter_1),
	.datac(!m0_write1),
	.datad(!uav_read),
	.datae(!av_waitrequest_generated),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_latency_shift_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~0 .extended_lut = "off";
defparam \read_latency_shift_reg~0 .lut_mask = 64'hDFFFFFFFDFFFFFFF;
defparam \read_latency_shift_reg~0 .shared_arith = "off";

endmodule

module first_nios2_system_altera_merlin_slave_translator_9 (
	av_readdata_pre_0,
	av_readdata_pre_1,
	av_readdata_pre_2,
	av_readdata_pre_3,
	av_readdata_pre_4,
	av_readdata_pre_5,
	av_readdata_pre_6,
	av_readdata_pre_7,
	av_readdata_pre_22,
	av_readdata_pre_21,
	av_readdata_pre_20,
	av_readdata_pre_19,
	av_readdata_pre_17,
	av_readdata_pre_18,
	av_readdata_pre_16,
	q_b_0,
	q_b_1,
	q_b_2,
	q_b_3,
	q_b_4,
	q_b_5,
	q_b_6,
	q_b_7,
	av_readdata,
	reset,
	read_latency_shift_reg,
	read_latency_shift_reg_0,
	av_waitrequest,
	av_waitrequest1,
	b_full,
	b_full1,
	read_0,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_5,
	av_readdata_pre_10,
	av_readdata_pre_8,
	av_readdata_pre_9,
	av_readdata_pre_15,
	av_readdata_pre_12,
	av_readdata_pre_13,
	av_readdata_pre_14,
	clk)/* synthesis synthesis_greybox=1 */;
output 	av_readdata_pre_0;
output 	av_readdata_pre_1;
output 	av_readdata_pre_2;
output 	av_readdata_pre_3;
output 	av_readdata_pre_4;
output 	av_readdata_pre_5;
output 	av_readdata_pre_6;
output 	av_readdata_pre_7;
output 	av_readdata_pre_22;
output 	av_readdata_pre_21;
output 	av_readdata_pre_20;
output 	av_readdata_pre_19;
output 	av_readdata_pre_17;
output 	av_readdata_pre_18;
output 	av_readdata_pre_16;
input 	q_b_0;
input 	q_b_1;
input 	q_b_2;
input 	q_b_3;
input 	q_b_4;
input 	q_b_5;
input 	q_b_6;
input 	q_b_7;
input 	[31:0] av_readdata;
input 	reset;
input 	read_latency_shift_reg;
output 	read_latency_shift_reg_0;
input 	av_waitrequest;
input 	av_waitrequest1;
input 	b_full;
input 	b_full1;
input 	read_0;
input 	counter_reg_bit_0;
input 	counter_reg_bit_1;
input 	counter_reg_bit_4;
input 	counter_reg_bit_3;
input 	counter_reg_bit_2;
input 	counter_reg_bit_5;
output 	av_readdata_pre_10;
output 	av_readdata_pre_8;
output 	av_readdata_pre_9;
output 	av_readdata_pre_15;
output 	av_readdata_pre_12;
output 	av_readdata_pre_13;
output 	av_readdata_pre_14;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read_latency_shift_reg~0_combout ;
wire \av_readdata_pre[13]~0_combout ;


dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(q_b_0),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

dffeas \av_readdata_pre[1] (
	.clk(clk),
	.d(av_readdata[1]),
	.asdata(q_b_1),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_1),
	.prn(vcc));
defparam \av_readdata_pre[1] .is_wysiwyg = "true";
defparam \av_readdata_pre[1] .power_up = "low";

dffeas \av_readdata_pre[2] (
	.clk(clk),
	.d(av_readdata[2]),
	.asdata(q_b_2),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_2),
	.prn(vcc));
defparam \av_readdata_pre[2] .is_wysiwyg = "true";
defparam \av_readdata_pre[2] .power_up = "low";

dffeas \av_readdata_pre[3] (
	.clk(clk),
	.d(av_readdata[2]),
	.asdata(q_b_3),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_3),
	.prn(vcc));
defparam \av_readdata_pre[3] .is_wysiwyg = "true";
defparam \av_readdata_pre[3] .power_up = "low";

dffeas \av_readdata_pre[4] (
	.clk(clk),
	.d(av_readdata[2]),
	.asdata(q_b_4),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_4),
	.prn(vcc));
defparam \av_readdata_pre[4] .is_wysiwyg = "true";
defparam \av_readdata_pre[4] .power_up = "low";

dffeas \av_readdata_pre[5] (
	.clk(clk),
	.d(av_readdata[2]),
	.asdata(q_b_5),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_5),
	.prn(vcc));
defparam \av_readdata_pre[5] .is_wysiwyg = "true";
defparam \av_readdata_pre[5] .power_up = "low";

dffeas \av_readdata_pre[6] (
	.clk(clk),
	.d(av_readdata[2]),
	.asdata(q_b_6),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_6),
	.prn(vcc));
defparam \av_readdata_pre[6] .is_wysiwyg = "true";
defparam \av_readdata_pre[6] .power_up = "low";

dffeas \av_readdata_pre[7] (
	.clk(clk),
	.d(av_readdata[2]),
	.asdata(q_b_7),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_7),
	.prn(vcc));
defparam \av_readdata_pre[7] .is_wysiwyg = "true";
defparam \av_readdata_pre[7] .power_up = "low";

dffeas \av_readdata_pre[22] (
	.clk(clk),
	.d(av_readdata[22]),
	.asdata(b_full),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_22),
	.prn(vcc));
defparam \av_readdata_pre[22] .is_wysiwyg = "true";
defparam \av_readdata_pre[22] .power_up = "low";

dffeas \av_readdata_pre[21] (
	.clk(clk),
	.d(av_readdata[21]),
	.asdata(counter_reg_bit_5),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_21),
	.prn(vcc));
defparam \av_readdata_pre[21] .is_wysiwyg = "true";
defparam \av_readdata_pre[21] .power_up = "low";

dffeas \av_readdata_pre[20] (
	.clk(clk),
	.d(av_readdata[20]),
	.asdata(counter_reg_bit_4),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_20),
	.prn(vcc));
defparam \av_readdata_pre[20] .is_wysiwyg = "true";
defparam \av_readdata_pre[20] .power_up = "low";

dffeas \av_readdata_pre[19] (
	.clk(clk),
	.d(av_readdata[19]),
	.asdata(counter_reg_bit_3),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_19),
	.prn(vcc));
defparam \av_readdata_pre[19] .is_wysiwyg = "true";
defparam \av_readdata_pre[19] .power_up = "low";

dffeas \av_readdata_pre[17] (
	.clk(clk),
	.d(av_readdata[17]),
	.asdata(counter_reg_bit_1),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_17),
	.prn(vcc));
defparam \av_readdata_pre[17] .is_wysiwyg = "true";
defparam \av_readdata_pre[17] .power_up = "low";

dffeas \av_readdata_pre[18] (
	.clk(clk),
	.d(av_readdata[18]),
	.asdata(counter_reg_bit_2),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_18),
	.prn(vcc));
defparam \av_readdata_pre[18] .is_wysiwyg = "true";
defparam \av_readdata_pre[18] .power_up = "low";

dffeas \av_readdata_pre[16] (
	.clk(clk),
	.d(av_readdata[16]),
	.asdata(counter_reg_bit_0),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_16),
	.prn(vcc));
defparam \av_readdata_pre[16] .is_wysiwyg = "true";
defparam \av_readdata_pre[16] .power_up = "low";

dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(\read_latency_shift_reg~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

dffeas \av_readdata_pre[10] (
	.clk(clk),
	.d(av_readdata[10]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_10),
	.prn(vcc));
defparam \av_readdata_pre[10] .is_wysiwyg = "true";
defparam \av_readdata_pre[10] .power_up = "low";

dffeas \av_readdata_pre[8] (
	.clk(clk),
	.d(av_readdata[8]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_8),
	.prn(vcc));
defparam \av_readdata_pre[8] .is_wysiwyg = "true";
defparam \av_readdata_pre[8] .power_up = "low";

dffeas \av_readdata_pre[9] (
	.clk(clk),
	.d(av_readdata[9]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_9),
	.prn(vcc));
defparam \av_readdata_pre[9] .is_wysiwyg = "true";
defparam \av_readdata_pre[9] .power_up = "low";

dffeas \av_readdata_pre[15] (
	.clk(clk),
	.d(av_readdata[15]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_15),
	.prn(vcc));
defparam \av_readdata_pre[15] .is_wysiwyg = "true";
defparam \av_readdata_pre[15] .power_up = "low";

dffeas \av_readdata_pre[12] (
	.clk(clk),
	.d(av_readdata[12]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_12),
	.prn(vcc));
defparam \av_readdata_pre[12] .is_wysiwyg = "true";
defparam \av_readdata_pre[12] .power_up = "low";

dffeas \av_readdata_pre[13] (
	.clk(clk),
	.d(\av_readdata_pre[13]~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_13),
	.prn(vcc));
defparam \av_readdata_pre[13] .is_wysiwyg = "true";
defparam \av_readdata_pre[13] .power_up = "low";

dffeas \av_readdata_pre[14] (
	.clk(clk),
	.d(av_readdata[14]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_14),
	.prn(vcc));
defparam \av_readdata_pre[14] .is_wysiwyg = "true";
defparam \av_readdata_pre[14] .power_up = "low";

cyclonev_lcell_comb \read_latency_shift_reg~0 (
	.dataa(!av_waitrequest),
	.datab(!av_waitrequest1),
	.datac(!read_latency_shift_reg),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_latency_shift_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~0 .extended_lut = "off";
defparam \read_latency_shift_reg~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \read_latency_shift_reg~0 .shared_arith = "off";

cyclonev_lcell_comb \av_readdata_pre[13]~0 (
	.dataa(!b_full1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_readdata_pre[13]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_readdata_pre[13]~0 .extended_lut = "off";
defparam \av_readdata_pre[13]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \av_readdata_pre[13]~0 .shared_arith = "off";

endmodule

module first_nios2_system_altera_merlin_slave_translator_10 (
	av_readdata_pre_0,
	av_readdata_pre_1,
	av_readdata_pre_2,
	av_readdata_pre_3,
	av_readdata_pre_4,
	av_readdata_pre_5,
	av_readdata_pre_6,
	av_readdata_pre_7,
	av_readdata,
	clr_break_line,
	d_write,
	Equal0,
	reset,
	wait_latency_counter_1,
	wait_latency_counter_0,
	m0_write,
	uav_read,
	cp_valid,
	read_latency_shift_reg_0,
	m0_write1,
	av_waitrequest_generated,
	clk)/* synthesis synthesis_greybox=1 */;
output 	av_readdata_pre_0;
output 	av_readdata_pre_1;
output 	av_readdata_pre_2;
output 	av_readdata_pre_3;
output 	av_readdata_pre_4;
output 	av_readdata_pre_5;
output 	av_readdata_pre_6;
output 	av_readdata_pre_7;
input 	[31:0] av_readdata;
input 	clr_break_line;
input 	d_write;
input 	Equal0;
input 	reset;
output 	wait_latency_counter_1;
output 	wait_latency_counter_0;
input 	m0_write;
input 	uav_read;
input 	cp_valid;
output 	read_latency_shift_reg_0;
input 	m0_write1;
output 	av_waitrequest_generated;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wait_latency_counter~0_combout ;
wire \wait_latency_counter~1_combout ;
wire \read_latency_shift_reg~0_combout ;


dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(Equal0),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

dffeas \av_readdata_pre[1] (
	.clk(clk),
	.d(av_readdata[1]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(Equal0),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_1),
	.prn(vcc));
defparam \av_readdata_pre[1] .is_wysiwyg = "true";
defparam \av_readdata_pre[1] .power_up = "low";

dffeas \av_readdata_pre[2] (
	.clk(clk),
	.d(av_readdata[2]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(Equal0),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_2),
	.prn(vcc));
defparam \av_readdata_pre[2] .is_wysiwyg = "true";
defparam \av_readdata_pre[2] .power_up = "low";

dffeas \av_readdata_pre[3] (
	.clk(clk),
	.d(av_readdata[3]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(Equal0),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_3),
	.prn(vcc));
defparam \av_readdata_pre[3] .is_wysiwyg = "true";
defparam \av_readdata_pre[3] .power_up = "low";

dffeas \av_readdata_pre[4] (
	.clk(clk),
	.d(av_readdata[4]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(Equal0),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_4),
	.prn(vcc));
defparam \av_readdata_pre[4] .is_wysiwyg = "true";
defparam \av_readdata_pre[4] .power_up = "low";

dffeas \av_readdata_pre[5] (
	.clk(clk),
	.d(av_readdata[5]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(Equal0),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_5),
	.prn(vcc));
defparam \av_readdata_pre[5] .is_wysiwyg = "true";
defparam \av_readdata_pre[5] .power_up = "low";

dffeas \av_readdata_pre[6] (
	.clk(clk),
	.d(av_readdata[6]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(Equal0),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_6),
	.prn(vcc));
defparam \av_readdata_pre[6] .is_wysiwyg = "true";
defparam \av_readdata_pre[6] .power_up = "low";

dffeas \av_readdata_pre[7] (
	.clk(clk),
	.d(av_readdata[7]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(Equal0),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_7),
	.prn(vcc));
defparam \av_readdata_pre[7] .is_wysiwyg = "true";
defparam \av_readdata_pre[7] .power_up = "low";

dffeas \wait_latency_counter[1] (
	.clk(clk),
	.d(\wait_latency_counter~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_1),
	.prn(vcc));
defparam \wait_latency_counter[1] .is_wysiwyg = "true";
defparam \wait_latency_counter[1] .power_up = "low";

dffeas \wait_latency_counter[0] (
	.clk(clk),
	.d(\wait_latency_counter~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_0),
	.prn(vcc));
defparam \wait_latency_counter[0] .is_wysiwyg = "true";
defparam \wait_latency_counter[0] .power_up = "low";

dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(\read_latency_shift_reg~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

cyclonev_lcell_comb \av_waitrequest_generated~0 (
	.dataa(!wait_latency_counter_0),
	.datab(!wait_latency_counter_1),
	.datac(!m0_write1),
	.datad(!m0_write),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(av_waitrequest_generated),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_waitrequest_generated~0 .extended_lut = "off";
defparam \av_waitrequest_generated~0 .lut_mask = 64'hEDDEEDDEEDDEEDDE;
defparam \av_waitrequest_generated~0 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter~0 (
	.dataa(!d_write),
	.datab(!wait_latency_counter_0),
	.datac(!wait_latency_counter_1),
	.datad(!m0_write1),
	.datae(!cp_valid),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~0 .extended_lut = "off";
defparam \wait_latency_counter~0 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \wait_latency_counter~0 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter~1 (
	.dataa(!wait_latency_counter_0),
	.datab(!m0_write1),
	.datac(!cp_valid),
	.datad(!av_waitrequest_generated),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~1 .extended_lut = "off";
defparam \wait_latency_counter~1 .lut_mask = 64'hFFBFFFBFFFBFFFBF;
defparam \wait_latency_counter~1 .shared_arith = "off";

cyclonev_lcell_comb \read_latency_shift_reg~0 (
	.dataa(!clr_break_line),
	.datab(!d_write),
	.datac(!wait_latency_counter_0),
	.datad(!wait_latency_counter_1),
	.datae(!m0_write1),
	.dataf(!uav_read),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_latency_shift_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~0 .extended_lut = "off";
defparam \read_latency_shift_reg~0 .lut_mask = 64'hFF7DFFFFFFFFFFFF;
defparam \read_latency_shift_reg~0 .shared_arith = "off";

endmodule

module first_nios2_system_altera_merlin_slave_translator_11 (
	clr_break_line,
	reset,
	read_latency_shift_reg_0,
	mem_used_1,
	WideOr1,
	mem,
	read_latency_shift_reg,
	clk)/* synthesis synthesis_greybox=1 */;
input 	clr_break_line;
input 	reset;
output 	read_latency_shift_reg_0;
input 	mem_used_1;
input 	WideOr1;
input 	mem;
output 	read_latency_shift_reg;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read_latency_shift_reg~1_combout ;


dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(\read_latency_shift_reg~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

cyclonev_lcell_comb \read_latency_shift_reg~0 (
	.dataa(!clr_break_line),
	.datab(!mem_used_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(read_latency_shift_reg),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~0 .extended_lut = "off";
defparam \read_latency_shift_reg~0 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \read_latency_shift_reg~0 .shared_arith = "off";

cyclonev_lcell_comb \read_latency_shift_reg~1 (
	.dataa(!WideOr1),
	.datab(!mem),
	.datac(!read_latency_shift_reg),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_latency_shift_reg~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~1 .extended_lut = "off";
defparam \read_latency_shift_reg~1 .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \read_latency_shift_reg~1 .shared_arith = "off";

endmodule

module first_nios2_system_altera_merlin_slave_translator_12 (
	av_readdata,
	d_write,
	reset,
	cp_valid,
	read_latency_shift_reg_0,
	wait_latency_counter_1,
	wait_latency_counter_0,
	sink_ready,
	m0_write,
	av_readdata_pre_0,
	clk)/* synthesis synthesis_greybox=1 */;
input 	[31:0] av_readdata;
input 	d_write;
input 	reset;
input 	cp_valid;
output 	read_latency_shift_reg_0;
output 	wait_latency_counter_1;
output 	wait_latency_counter_0;
input 	sink_ready;
input 	m0_write;
output 	av_readdata_pre_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wait_latency_counter~0_combout ;
wire \wait_latency_counter~1_combout ;


dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(sink_ready),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

dffeas \wait_latency_counter[1] (
	.clk(clk),
	.d(\wait_latency_counter~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_1),
	.prn(vcc));
defparam \wait_latency_counter[1] .is_wysiwyg = "true";
defparam \wait_latency_counter[1] .power_up = "low";

dffeas \wait_latency_counter[0] (
	.clk(clk),
	.d(\wait_latency_counter~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_0),
	.prn(vcc));
defparam \wait_latency_counter[0] .is_wysiwyg = "true";
defparam \wait_latency_counter[0] .power_up = "low";

dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

cyclonev_lcell_comb \wait_latency_counter~0 (
	.dataa(!d_write),
	.datab(!cp_valid),
	.datac(!wait_latency_counter_1),
	.datad(!wait_latency_counter_0),
	.datae(!m0_write),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~0 .extended_lut = "off";
defparam \wait_latency_counter~0 .lut_mask = 64'h7FF7FFFF7FF7FFFF;
defparam \wait_latency_counter~0 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter~1 (
	.dataa(!d_write),
	.datab(!cp_valid),
	.datac(!wait_latency_counter_1),
	.datad(!wait_latency_counter_0),
	.datae(!m0_write),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~1 .extended_lut = "off";
defparam \wait_latency_counter~1 .lut_mask = 64'hFFBFFFFFFFBFFFFF;
defparam \wait_latency_counter~1 .shared_arith = "off";

endmodule

module first_nios2_system_altera_merlin_slave_translator_13 (
	av_readdata,
	d_write,
	reset,
	cp_valid,
	read_latency_shift_reg_0,
	wait_latency_counter_1,
	wait_latency_counter_0,
	sink_ready,
	m0_write,
	av_readdata_pre_0,
	clk)/* synthesis synthesis_greybox=1 */;
input 	[31:0] av_readdata;
input 	d_write;
input 	reset;
input 	cp_valid;
output 	read_latency_shift_reg_0;
output 	wait_latency_counter_1;
output 	wait_latency_counter_0;
input 	sink_ready;
input 	m0_write;
output 	av_readdata_pre_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wait_latency_counter~0_combout ;
wire \wait_latency_counter~1_combout ;


dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(sink_ready),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

dffeas \wait_latency_counter[1] (
	.clk(clk),
	.d(\wait_latency_counter~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_1),
	.prn(vcc));
defparam \wait_latency_counter[1] .is_wysiwyg = "true";
defparam \wait_latency_counter[1] .power_up = "low";

dffeas \wait_latency_counter[0] (
	.clk(clk),
	.d(\wait_latency_counter~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_0),
	.prn(vcc));
defparam \wait_latency_counter[0] .is_wysiwyg = "true";
defparam \wait_latency_counter[0] .power_up = "low";

dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

cyclonev_lcell_comb \wait_latency_counter~0 (
	.dataa(!d_write),
	.datab(!cp_valid),
	.datac(!wait_latency_counter_1),
	.datad(!wait_latency_counter_0),
	.datae(!m0_write),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~0 .extended_lut = "off";
defparam \wait_latency_counter~0 .lut_mask = 64'h7FF7FFFF7FF7FFFF;
defparam \wait_latency_counter~0 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter~1 (
	.dataa(!d_write),
	.datab(!cp_valid),
	.datac(!wait_latency_counter_1),
	.datad(!wait_latency_counter_0),
	.datae(!m0_write),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~1 .extended_lut = "off";
defparam \wait_latency_counter~1 .lut_mask = 64'hFFBFFFFFFFBFFFFF;
defparam \wait_latency_counter~1 .shared_arith = "off";

endmodule

module first_nios2_system_altera_merlin_slave_translator_14 (
	av_readdata_pre_0,
	av_readdata,
	clr_break_line,
	d_write,
	Equal0,
	reset,
	wait_latency_counter_1,
	m0_write,
	wait_latency_counter_0,
	m0_write1,
	uav_read,
	cp_valid,
	read_latency_shift_reg_0,
	av_waitrequest_generated,
	clk)/* synthesis synthesis_greybox=1 */;
output 	av_readdata_pre_0;
input 	[31:0] av_readdata;
input 	clr_break_line;
input 	d_write;
input 	Equal0;
input 	reset;
output 	wait_latency_counter_1;
input 	m0_write;
output 	wait_latency_counter_0;
input 	m0_write1;
input 	uav_read;
input 	cp_valid;
output 	read_latency_shift_reg_0;
output 	av_waitrequest_generated;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wait_latency_counter~0_combout ;
wire \wait_latency_counter~1_combout ;
wire \read_latency_shift_reg~0_combout ;


dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(Equal0),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

dffeas \wait_latency_counter[1] (
	.clk(clk),
	.d(\wait_latency_counter~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_1),
	.prn(vcc));
defparam \wait_latency_counter[1] .is_wysiwyg = "true";
defparam \wait_latency_counter[1] .power_up = "low";

dffeas \wait_latency_counter[0] (
	.clk(clk),
	.d(\wait_latency_counter~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_0),
	.prn(vcc));
defparam \wait_latency_counter[0] .is_wysiwyg = "true";
defparam \wait_latency_counter[0] .power_up = "low";

dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(\read_latency_shift_reg~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

cyclonev_lcell_comb \av_waitrequest_generated~0 (
	.dataa(!wait_latency_counter_0),
	.datab(!wait_latency_counter_1),
	.datac(!m0_write),
	.datad(!m0_write1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(av_waitrequest_generated),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_waitrequest_generated~0 .extended_lut = "off";
defparam \av_waitrequest_generated~0 .lut_mask = 64'hEDDEEDDEEDDEEDDE;
defparam \av_waitrequest_generated~0 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter~0 (
	.dataa(!d_write),
	.datab(!wait_latency_counter_0),
	.datac(!wait_latency_counter_1),
	.datad(!m0_write),
	.datae(!cp_valid),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~0 .extended_lut = "off";
defparam \wait_latency_counter~0 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \wait_latency_counter~0 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter~1 (
	.dataa(!wait_latency_counter_0),
	.datab(!m0_write),
	.datac(!cp_valid),
	.datad(!av_waitrequest_generated),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~1 .extended_lut = "off";
defparam \wait_latency_counter~1 .lut_mask = 64'hFFBFFFBFFFBFFFBF;
defparam \wait_latency_counter~1 .shared_arith = "off";

cyclonev_lcell_comb \read_latency_shift_reg~0 (
	.dataa(!clr_break_line),
	.datab(!d_write),
	.datac(!wait_latency_counter_0),
	.datad(!wait_latency_counter_1),
	.datae(!m0_write),
	.dataf(!uav_read),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_latency_shift_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~0 .extended_lut = "off";
defparam \read_latency_shift_reg~0 .lut_mask = 64'hFF7DFFFFFFFFFFFF;
defparam \read_latency_shift_reg~0 .shared_arith = "off";

endmodule

module first_nios2_system_altera_merlin_slave_translator_15 (
	clr_break_line,
	d_write,
	reset,
	m0_write,
	uav_read,
	cp_valid,
	read_latency_shift_reg_0,
	wait_latency_counter_0,
	wait_latency_counter_1,
	m0_write1,
	av_waitrequest_generated,
	av_readdata_pre_0,
	av_readdata_pre_1,
	av_readdata_pre_2,
	av_readdata_pre_3,
	av_readdata_pre_4,
	av_readdata_pre_5,
	av_readdata_pre_6,
	av_readdata_pre_7,
	av_readdata_pre_11,
	av_readdata_pre_10,
	av_readdata_pre_8,
	av_readdata_pre_9,
	av_readdata_pre_15,
	av_readdata_pre_12,
	av_readdata_pre_13,
	av_readdata_pre_14,
	av_readdata,
	clk)/* synthesis synthesis_greybox=1 */;
input 	clr_break_line;
input 	d_write;
input 	reset;
input 	m0_write;
input 	uav_read;
input 	cp_valid;
output 	read_latency_shift_reg_0;
output 	wait_latency_counter_0;
output 	wait_latency_counter_1;
input 	m0_write1;
output 	av_waitrequest_generated;
output 	av_readdata_pre_0;
output 	av_readdata_pre_1;
output 	av_readdata_pre_2;
output 	av_readdata_pre_3;
output 	av_readdata_pre_4;
output 	av_readdata_pre_5;
output 	av_readdata_pre_6;
output 	av_readdata_pre_7;
output 	av_readdata_pre_11;
output 	av_readdata_pre_10;
output 	av_readdata_pre_8;
output 	av_readdata_pre_9;
output 	av_readdata_pre_15;
output 	av_readdata_pre_12;
output 	av_readdata_pre_13;
output 	av_readdata_pre_14;
input 	[31:0] av_readdata;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read_latency_shift_reg~0_combout ;
wire \wait_latency_counter~0_combout ;
wire \wait_latency_counter~1_combout ;


dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(\read_latency_shift_reg~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

dffeas \wait_latency_counter[0] (
	.clk(clk),
	.d(\wait_latency_counter~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_0),
	.prn(vcc));
defparam \wait_latency_counter[0] .is_wysiwyg = "true";
defparam \wait_latency_counter[0] .power_up = "low";

dffeas \wait_latency_counter[1] (
	.clk(clk),
	.d(\wait_latency_counter~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_1),
	.prn(vcc));
defparam \wait_latency_counter[1] .is_wysiwyg = "true";
defparam \wait_latency_counter[1] .power_up = "low";

cyclonev_lcell_comb \av_waitrequest_generated~0 (
	.dataa(!m0_write),
	.datab(!wait_latency_counter_0),
	.datac(!m0_write1),
	.datad(!wait_latency_counter_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(av_waitrequest_generated),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_waitrequest_generated~0 .extended_lut = "off";
defparam \av_waitrequest_generated~0 .lut_mask = 64'hFF96FF96FF96FF96;
defparam \av_waitrequest_generated~0 .shared_arith = "off";

dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

dffeas \av_readdata_pre[1] (
	.clk(clk),
	.d(av_readdata[1]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_1),
	.prn(vcc));
defparam \av_readdata_pre[1] .is_wysiwyg = "true";
defparam \av_readdata_pre[1] .power_up = "low";

dffeas \av_readdata_pre[2] (
	.clk(clk),
	.d(av_readdata[2]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_2),
	.prn(vcc));
defparam \av_readdata_pre[2] .is_wysiwyg = "true";
defparam \av_readdata_pre[2] .power_up = "low";

dffeas \av_readdata_pre[3] (
	.clk(clk),
	.d(av_readdata[3]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_3),
	.prn(vcc));
defparam \av_readdata_pre[3] .is_wysiwyg = "true";
defparam \av_readdata_pre[3] .power_up = "low";

dffeas \av_readdata_pre[4] (
	.clk(clk),
	.d(av_readdata[4]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_4),
	.prn(vcc));
defparam \av_readdata_pre[4] .is_wysiwyg = "true";
defparam \av_readdata_pre[4] .power_up = "low";

dffeas \av_readdata_pre[5] (
	.clk(clk),
	.d(av_readdata[5]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_5),
	.prn(vcc));
defparam \av_readdata_pre[5] .is_wysiwyg = "true";
defparam \av_readdata_pre[5] .power_up = "low";

dffeas \av_readdata_pre[6] (
	.clk(clk),
	.d(av_readdata[6]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_6),
	.prn(vcc));
defparam \av_readdata_pre[6] .is_wysiwyg = "true";
defparam \av_readdata_pre[6] .power_up = "low";

dffeas \av_readdata_pre[7] (
	.clk(clk),
	.d(av_readdata[7]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_7),
	.prn(vcc));
defparam \av_readdata_pre[7] .is_wysiwyg = "true";
defparam \av_readdata_pre[7] .power_up = "low";

dffeas \av_readdata_pre[11] (
	.clk(clk),
	.d(av_readdata[11]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_11),
	.prn(vcc));
defparam \av_readdata_pre[11] .is_wysiwyg = "true";
defparam \av_readdata_pre[11] .power_up = "low";

dffeas \av_readdata_pre[10] (
	.clk(clk),
	.d(av_readdata[10]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_10),
	.prn(vcc));
defparam \av_readdata_pre[10] .is_wysiwyg = "true";
defparam \av_readdata_pre[10] .power_up = "low";

dffeas \av_readdata_pre[8] (
	.clk(clk),
	.d(av_readdata[8]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_8),
	.prn(vcc));
defparam \av_readdata_pre[8] .is_wysiwyg = "true";
defparam \av_readdata_pre[8] .power_up = "low";

dffeas \av_readdata_pre[9] (
	.clk(clk),
	.d(av_readdata[9]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_9),
	.prn(vcc));
defparam \av_readdata_pre[9] .is_wysiwyg = "true";
defparam \av_readdata_pre[9] .power_up = "low";

dffeas \av_readdata_pre[15] (
	.clk(clk),
	.d(av_readdata[15]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_15),
	.prn(vcc));
defparam \av_readdata_pre[15] .is_wysiwyg = "true";
defparam \av_readdata_pre[15] .power_up = "low";

dffeas \av_readdata_pre[12] (
	.clk(clk),
	.d(av_readdata[12]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_12),
	.prn(vcc));
defparam \av_readdata_pre[12] .is_wysiwyg = "true";
defparam \av_readdata_pre[12] .power_up = "low";

dffeas \av_readdata_pre[13] (
	.clk(clk),
	.d(av_readdata[13]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_13),
	.prn(vcc));
defparam \av_readdata_pre[13] .is_wysiwyg = "true";
defparam \av_readdata_pre[13] .power_up = "low";

dffeas \av_readdata_pre[14] (
	.clk(clk),
	.d(av_readdata[14]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_14),
	.prn(vcc));
defparam \av_readdata_pre[14] .is_wysiwyg = "true";
defparam \av_readdata_pre[14] .power_up = "low";

cyclonev_lcell_comb \read_latency_shift_reg~0 (
	.dataa(!clr_break_line),
	.datab(!d_write),
	.datac(!uav_read),
	.datad(!wait_latency_counter_0),
	.datae(!m0_write1),
	.dataf(!wait_latency_counter_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_latency_shift_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~0 .extended_lut = "off";
defparam \read_latency_shift_reg~0 .lut_mask = 64'hFFFFFFFF7FDFFFFF;
defparam \read_latency_shift_reg~0 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter~0 (
	.dataa(!cp_valid),
	.datab(!wait_latency_counter_0),
	.datac(!m0_write1),
	.datad(!av_waitrequest_generated),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~0 .extended_lut = "off";
defparam \wait_latency_counter~0 .lut_mask = 64'hFFDFFFDFFFDFFFDF;
defparam \wait_latency_counter~0 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter~1 (
	.dataa(!d_write),
	.datab(!cp_valid),
	.datac(!wait_latency_counter_0),
	.datad(!m0_write1),
	.datae(!wait_latency_counter_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~1 .extended_lut = "off";
defparam \wait_latency_counter~1 .lut_mask = 64'h7FFFF7FF7FFFF7FF;
defparam \wait_latency_counter~1 .shared_arith = "off";

endmodule

module first_nios2_system_altera_merlin_slave_translator_16 (
	d_write,
	av_readdata,
	reset,
	cp_valid,
	read_latency_shift_reg_0,
	mem_used_1,
	wait_latency_counter_1,
	wait_latency_counter_0,
	always1,
	sink_ready,
	av_readdata_pre_30,
	clk)/* synthesis synthesis_greybox=1 */;
input 	d_write;
input 	[31:0] av_readdata;
input 	reset;
input 	cp_valid;
output 	read_latency_shift_reg_0;
input 	mem_used_1;
output 	wait_latency_counter_1;
output 	wait_latency_counter_0;
input 	always1;
input 	sink_ready;
output 	av_readdata_pre_30;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wait_latency_counter[1]~0_combout ;
wire \wait_latency_counter~1_combout ;
wire \wait_latency_counter~2_combout ;


dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(sink_ready),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

dffeas \wait_latency_counter[1] (
	.clk(clk),
	.d(\wait_latency_counter~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_1),
	.prn(vcc));
defparam \wait_latency_counter[1] .is_wysiwyg = "true";
defparam \wait_latency_counter[1] .power_up = "low";

dffeas \wait_latency_counter[0] (
	.clk(clk),
	.d(\wait_latency_counter~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_0),
	.prn(vcc));
defparam \wait_latency_counter[0] .is_wysiwyg = "true";
defparam \wait_latency_counter[0] .power_up = "low";

dffeas \av_readdata_pre[30] (
	.clk(clk),
	.d(av_readdata[30]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_30),
	.prn(vcc));
defparam \av_readdata_pre[30] .is_wysiwyg = "true";
defparam \av_readdata_pre[30] .power_up = "low";

cyclonev_lcell_comb \wait_latency_counter[1]~0 (
	.dataa(!d_write),
	.datab(!cp_valid),
	.datac(!mem_used_1),
	.datad(!wait_latency_counter_1),
	.datae(!wait_latency_counter_0),
	.dataf(!always1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter[1]~0 .extended_lut = "off";
defparam \wait_latency_counter[1]~0 .lut_mask = 64'hF7FFFBFFFFFFFFFF;
defparam \wait_latency_counter[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter~1 (
	.dataa(!wait_latency_counter_1),
	.datab(!wait_latency_counter_0),
	.datac(!\wait_latency_counter[1]~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~1 .extended_lut = "off";
defparam \wait_latency_counter~1 .lut_mask = 64'h6F6F6F6F6F6F6F6F;
defparam \wait_latency_counter~1 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter~2 (
	.dataa(!wait_latency_counter_0),
	.datab(!\wait_latency_counter[1]~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~2 .extended_lut = "off";
defparam \wait_latency_counter~2 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \wait_latency_counter~2 .shared_arith = "off";

endmodule

module first_nios2_system_altera_merlin_slave_translator_17 (
	av_readdata,
	d_write,
	reset,
	cp_valid,
	read_latency_shift_reg_0,
	wait_latency_counter_1,
	wait_latency_counter_0,
	sink_ready,
	m0_write,
	av_readdata_pre_0,
	av_readdata_pre_1,
	av_readdata_pre_2,
	av_readdata_pre_3,
	clk)/* synthesis synthesis_greybox=1 */;
input 	[31:0] av_readdata;
input 	d_write;
input 	reset;
input 	cp_valid;
output 	read_latency_shift_reg_0;
output 	wait_latency_counter_1;
output 	wait_latency_counter_0;
input 	sink_ready;
input 	m0_write;
output 	av_readdata_pre_0;
output 	av_readdata_pre_1;
output 	av_readdata_pre_2;
output 	av_readdata_pre_3;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wait_latency_counter~0_combout ;
wire \wait_latency_counter~1_combout ;


dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(sink_ready),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

dffeas \wait_latency_counter[1] (
	.clk(clk),
	.d(\wait_latency_counter~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_1),
	.prn(vcc));
defparam \wait_latency_counter[1] .is_wysiwyg = "true";
defparam \wait_latency_counter[1] .power_up = "low";

dffeas \wait_latency_counter[0] (
	.clk(clk),
	.d(\wait_latency_counter~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_0),
	.prn(vcc));
defparam \wait_latency_counter[0] .is_wysiwyg = "true";
defparam \wait_latency_counter[0] .power_up = "low";

dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

dffeas \av_readdata_pre[1] (
	.clk(clk),
	.d(av_readdata[1]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_1),
	.prn(vcc));
defparam \av_readdata_pre[1] .is_wysiwyg = "true";
defparam \av_readdata_pre[1] .power_up = "low";

dffeas \av_readdata_pre[2] (
	.clk(clk),
	.d(av_readdata[2]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_2),
	.prn(vcc));
defparam \av_readdata_pre[2] .is_wysiwyg = "true";
defparam \av_readdata_pre[2] .power_up = "low";

dffeas \av_readdata_pre[3] (
	.clk(clk),
	.d(av_readdata[3]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_3),
	.prn(vcc));
defparam \av_readdata_pre[3] .is_wysiwyg = "true";
defparam \av_readdata_pre[3] .power_up = "low";

cyclonev_lcell_comb \wait_latency_counter~0 (
	.dataa(!d_write),
	.datab(!cp_valid),
	.datac(!wait_latency_counter_1),
	.datad(!wait_latency_counter_0),
	.datae(!m0_write),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~0 .extended_lut = "off";
defparam \wait_latency_counter~0 .lut_mask = 64'h7FF7FFFF7FF7FFFF;
defparam \wait_latency_counter~0 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter~1 (
	.dataa(!d_write),
	.datab(!cp_valid),
	.datac(!wait_latency_counter_1),
	.datad(!wait_latency_counter_0),
	.datae(!m0_write),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~1 .extended_lut = "off";
defparam \wait_latency_counter~1 .lut_mask = 64'hFFBFFFFFFFBFFFFF;
defparam \wait_latency_counter~1 .shared_arith = "off";

endmodule

module first_nios2_system_altera_merlin_slave_translator_18 (
	av_readdata,
	d_write,
	reset,
	cp_valid,
	read_latency_shift_reg_0,
	wait_latency_counter_1,
	wait_latency_counter_0,
	sink_ready,
	m0_write,
	av_readdata_pre_0,
	av_readdata_pre_1,
	av_readdata_pre_2,
	av_readdata_pre_3,
	clk)/* synthesis synthesis_greybox=1 */;
input 	[31:0] av_readdata;
input 	d_write;
input 	reset;
input 	cp_valid;
output 	read_latency_shift_reg_0;
output 	wait_latency_counter_1;
output 	wait_latency_counter_0;
input 	sink_ready;
input 	m0_write;
output 	av_readdata_pre_0;
output 	av_readdata_pre_1;
output 	av_readdata_pre_2;
output 	av_readdata_pre_3;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wait_latency_counter~0_combout ;
wire \wait_latency_counter~1_combout ;


dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(sink_ready),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

dffeas \wait_latency_counter[1] (
	.clk(clk),
	.d(\wait_latency_counter~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_1),
	.prn(vcc));
defparam \wait_latency_counter[1] .is_wysiwyg = "true";
defparam \wait_latency_counter[1] .power_up = "low";

dffeas \wait_latency_counter[0] (
	.clk(clk),
	.d(\wait_latency_counter~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_0),
	.prn(vcc));
defparam \wait_latency_counter[0] .is_wysiwyg = "true";
defparam \wait_latency_counter[0] .power_up = "low";

dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

dffeas \av_readdata_pre[1] (
	.clk(clk),
	.d(av_readdata[1]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_1),
	.prn(vcc));
defparam \av_readdata_pre[1] .is_wysiwyg = "true";
defparam \av_readdata_pre[1] .power_up = "low";

dffeas \av_readdata_pre[2] (
	.clk(clk),
	.d(av_readdata[2]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_2),
	.prn(vcc));
defparam \av_readdata_pre[2] .is_wysiwyg = "true";
defparam \av_readdata_pre[2] .power_up = "low";

dffeas \av_readdata_pre[3] (
	.clk(clk),
	.d(av_readdata[3]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_3),
	.prn(vcc));
defparam \av_readdata_pre[3] .is_wysiwyg = "true";
defparam \av_readdata_pre[3] .power_up = "low";

cyclonev_lcell_comb \wait_latency_counter~0 (
	.dataa(!d_write),
	.datab(!cp_valid),
	.datac(!wait_latency_counter_1),
	.datad(!wait_latency_counter_0),
	.datae(!m0_write),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~0 .extended_lut = "off";
defparam \wait_latency_counter~0 .lut_mask = 64'h7FF7FFFF7FF7FFFF;
defparam \wait_latency_counter~0 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter~1 (
	.dataa(!d_write),
	.datab(!cp_valid),
	.datac(!wait_latency_counter_1),
	.datad(!wait_latency_counter_0),
	.datae(!m0_write),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~1 .extended_lut = "off";
defparam \wait_latency_counter~1 .lut_mask = 64'hFFBFFFFFFFBFFFFF;
defparam \wait_latency_counter~1 .shared_arith = "off";

endmodule

module first_nios2_system_altera_merlin_traffic_limiter (
	clr_break_line,
	reset,
	last_dest_id_2,
	has_pending_responses1,
	i_read,
	cmd_sink_data,
	last_dest_id_3,
	save_dest_id,
	WideOr0,
	nonposted_cmd_accepted1,
	src1_valid,
	src1_valid1,
	mem_61_0,
	mem_61_01,
	suppress_change_dest_id,
	clk)/* synthesis synthesis_greybox=1 */;
input 	clr_break_line;
input 	reset;
output 	last_dest_id_2;
output 	has_pending_responses1;
input 	i_read;
input 	[96:0] cmd_sink_data;
output 	last_dest_id_3;
output 	save_dest_id;
input 	WideOr0;
output 	nonposted_cmd_accepted1;
input 	src1_valid;
input 	src1_valid1;
input 	mem_61_0;
input 	mem_61_01;
output 	suppress_change_dest_id;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \response_sink_accepted~0_combout ;
wire \pending_response_count[0]~0_combout ;
wire \pending_response_count[0]~q ;
wire \has_pending_responses~0_combout ;
wire \last_dest_id[3]~0_combout ;


dffeas \last_dest_id[2] (
	.clk(clk),
	.d(cmd_sink_data[81]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(save_dest_id),
	.q(last_dest_id_2),
	.prn(vcc));
defparam \last_dest_id[2] .is_wysiwyg = "true";
defparam \last_dest_id[2] .power_up = "low";

dffeas has_pending_responses(
	.clk(clk),
	.d(\has_pending_responses~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(has_pending_responses1),
	.prn(vcc));
defparam has_pending_responses.is_wysiwyg = "true";
defparam has_pending_responses.power_up = "low";

dffeas \last_dest_id[3] (
	.clk(clk),
	.d(\last_dest_id[3]~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(save_dest_id),
	.q(last_dest_id_3),
	.prn(vcc));
defparam \last_dest_id[3] .is_wysiwyg = "true";
defparam \last_dest_id[3] .power_up = "low";

cyclonev_lcell_comb \save_dest_id~0 (
	.dataa(!clr_break_line),
	.datab(!last_dest_id_2),
	.datac(!has_pending_responses1),
	.datad(!i_read),
	.datae(!cmd_sink_data[81]),
	.dataf(!last_dest_id_3),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(save_dest_id),
	.sumout(),
	.cout(),
	.shareout());
defparam \save_dest_id~0 .extended_lut = "off";
defparam \save_dest_id~0 .lut_mask = 64'hFDFFF7FFF7FFFDFF;
defparam \save_dest_id~0 .shared_arith = "off";

cyclonev_lcell_comb nonposted_cmd_accepted(
	.dataa(!save_dest_id),
	.datab(!WideOr0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nonposted_cmd_accepted1),
	.sumout(),
	.cout(),
	.shareout());
defparam nonposted_cmd_accepted.extended_lut = "off";
defparam nonposted_cmd_accepted.lut_mask = 64'h7777777777777777;
defparam nonposted_cmd_accepted.shared_arith = "off";

cyclonev_lcell_comb \suppress_change_dest_id~0 (
	.dataa(!last_dest_id_2),
	.datab(!has_pending_responses1),
	.datac(!cmd_sink_data[81]),
	.datad(!last_dest_id_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(suppress_change_dest_id),
	.sumout(),
	.cout(),
	.shareout());
defparam \suppress_change_dest_id~0 .extended_lut = "off";
defparam \suppress_change_dest_id~0 .lut_mask = 64'hB77BB77BB77BB77B;
defparam \suppress_change_dest_id~0 .shared_arith = "off";

cyclonev_lcell_comb \response_sink_accepted~0 (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!mem_61_0),
	.datad(!mem_61_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\response_sink_accepted~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \response_sink_accepted~0 .extended_lut = "off";
defparam \response_sink_accepted~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \response_sink_accepted~0 .shared_arith = "off";

cyclonev_lcell_comb \pending_response_count[0]~0 (
	.dataa(!nonposted_cmd_accepted1),
	.datab(!\pending_response_count[0]~q ),
	.datac(!\response_sink_accepted~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pending_response_count[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pending_response_count[0]~0 .extended_lut = "off";
defparam \pending_response_count[0]~0 .lut_mask = 64'h9696969696969696;
defparam \pending_response_count[0]~0 .shared_arith = "off";

dffeas \pending_response_count[0] (
	.clk(clk),
	.d(\pending_response_count[0]~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\pending_response_count[0]~q ),
	.prn(vcc));
defparam \pending_response_count[0] .is_wysiwyg = "true";
defparam \pending_response_count[0] .power_up = "low";

cyclonev_lcell_comb \has_pending_responses~0 (
	.dataa(!has_pending_responses1),
	.datab(!nonposted_cmd_accepted1),
	.datac(!\pending_response_count[0]~q ),
	.datad(!\response_sink_accepted~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\has_pending_responses~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \has_pending_responses~0 .extended_lut = "off";
defparam \has_pending_responses~0 .lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam \has_pending_responses~0 .shared_arith = "off";

cyclonev_lcell_comb \last_dest_id[3]~0 (
	.dataa(!cmd_sink_data[81]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\last_dest_id[3]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_dest_id[3]~0 .extended_lut = "off";
defparam \last_dest_id[3]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \last_dest_id[3]~0 .shared_arith = "off";

endmodule

module first_nios2_system_first_nios2_system_mm_interconnect_0_cmd_demux (
	clr_break_line,
	wait_latency_counter_1,
	m0_write,
	wait_latency_counter_0,
	Equal6,
	wait_latency_counter_11,
	m0_write1,
	wait_latency_counter_01,
	m0_write2,
	cp_valid,
	write,
	write1,
	write2,
	mem_used_1,
	saved_grant_0,
	always1,
	src_channel_2,
	src_channel_21,
	Equal1,
	write3,
	write4,
	WideOr0,
	mem_used_11,
	wait_latency_counter_12,
	wait_latency_counter_02,
	always11,
	sink_ready,
	always12,
	mem_used_12,
	wait_latency_counter_13,
	wait_latency_counter_03,
	sink_ready1,
	always13,
	mem_used_13,
	wait_latency_counter_14,
	wait_latency_counter_04,
	sink_ready2,
	mem_used_14,
	av_waitrequest_generated,
	sink_ready3,
	mem_used_15,
	always14,
	av_waitrequest_generated1,
	sink_ready4,
	av_waitrequest,
	av_waitrequest1,
	mem_used_16,
	wait_latency_counter_15,
	wait_latency_counter_05,
	always15,
	sink_ready5,
	always16,
	mem_used_17,
	wait_latency_counter_16,
	wait_latency_counter_06,
	sink_ready6,
	mem_used_18,
	wait_latency_counter_17,
	wait_latency_counter_07,
	always17,
	sink_ready7,
	mem_used_19,
	wait_latency_counter_18,
	wait_latency_counter_08,
	always18,
	sink_ready8,
	saved_grant_01,
	write5,
	WideOr01,
	sink_ready9,
	sink_ready10,
	src3_valid,
	sink_ready11,
	sink_ready12,
	sink_ready13,
	sink_ready14,
	sink_ready15,
	sink_ready16,
	sink_ready17,
	src2_valid)/* synthesis synthesis_greybox=1 */;
input 	clr_break_line;
input 	wait_latency_counter_1;
input 	m0_write;
input 	wait_latency_counter_0;
input 	Equal6;
input 	wait_latency_counter_11;
input 	m0_write1;
input 	wait_latency_counter_01;
input 	m0_write2;
input 	cp_valid;
input 	write;
input 	write1;
input 	write2;
input 	mem_used_1;
input 	saved_grant_0;
input 	always1;
input 	src_channel_2;
input 	src_channel_21;
input 	Equal1;
input 	write3;
input 	write4;
output 	WideOr0;
input 	mem_used_11;
input 	wait_latency_counter_12;
input 	wait_latency_counter_02;
input 	always11;
output 	sink_ready;
input 	always12;
input 	mem_used_12;
input 	wait_latency_counter_13;
input 	wait_latency_counter_03;
output 	sink_ready1;
input 	always13;
input 	mem_used_13;
input 	wait_latency_counter_14;
input 	wait_latency_counter_04;
output 	sink_ready2;
input 	mem_used_14;
input 	av_waitrequest_generated;
output 	sink_ready3;
input 	mem_used_15;
input 	always14;
input 	av_waitrequest_generated1;
output 	sink_ready4;
input 	av_waitrequest;
input 	av_waitrequest1;
input 	mem_used_16;
input 	wait_latency_counter_15;
input 	wait_latency_counter_05;
input 	always15;
output 	sink_ready5;
input 	always16;
input 	mem_used_17;
input 	wait_latency_counter_16;
input 	wait_latency_counter_06;
output 	sink_ready6;
input 	mem_used_18;
input 	wait_latency_counter_17;
input 	wait_latency_counter_07;
input 	always17;
output 	sink_ready7;
input 	mem_used_19;
input 	wait_latency_counter_18;
input 	wait_latency_counter_08;
input 	always18;
output 	sink_ready8;
input 	saved_grant_01;
input 	write5;
output 	WideOr01;
output 	sink_ready9;
output 	sink_ready10;
output 	src3_valid;
output 	sink_ready11;
output 	sink_ready12;
output 	sink_ready13;
output 	sink_ready14;
output 	sink_ready15;
output 	sink_ready16;
output 	sink_ready17;
output 	src2_valid;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \WideOr0~0_combout ;
wire \WideOr0~1_combout ;
wire \WideOr0~2_combout ;
wire \WideOr0~4_combout ;
wire \WideOr0~5_combout ;
wire \sink_ready~9_combout ;


cyclonev_lcell_comb \WideOr0~3 (
	.dataa(!\WideOr0~0_combout ),
	.datab(!write),
	.datac(!write1),
	.datad(!write2),
	.datae(!\WideOr0~1_combout ),
	.dataf(!\WideOr0~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr0),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~3 .extended_lut = "off";
defparam \WideOr0~3 .lut_mask = 64'hFFFFFFFEFFFFFFFF;
defparam \WideOr0~3 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~0 (
	.dataa(!clr_break_line),
	.datab(!m0_write2),
	.datac(!mem_used_11),
	.datad(!wait_latency_counter_12),
	.datae(!wait_latency_counter_02),
	.dataf(!always11),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(sink_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~0 .extended_lut = "off";
defparam \sink_ready~0 .lut_mask = 64'hFFF7FFFDFFFFFFFF;
defparam \sink_ready~0 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~1 (
	.dataa(!clr_break_line),
	.datab(!m0_write2),
	.datac(!always12),
	.datad(!mem_used_12),
	.datae(!wait_latency_counter_13),
	.dataf(!wait_latency_counter_03),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(sink_ready1),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~1 .extended_lut = "off";
defparam \sink_ready~1 .lut_mask = 64'hFFFFFF7FFFFFFFDF;
defparam \sink_ready~1 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~2 (
	.dataa(!clr_break_line),
	.datab(!m0_write2),
	.datac(!always13),
	.datad(!mem_used_13),
	.datae(!wait_latency_counter_14),
	.dataf(!wait_latency_counter_04),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(sink_ready2),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~2 .extended_lut = "off";
defparam \sink_ready~2 .lut_mask = 64'hFFFFFF7FFFFFFFDF;
defparam \sink_ready~2 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~3 (
	.dataa(!clr_break_line),
	.datab(!Equal6),
	.datac(!always1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(sink_ready3),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~3 .extended_lut = "off";
defparam \sink_ready~3 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \sink_ready~3 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~4 (
	.dataa(!clr_break_line),
	.datab(!always1),
	.datac(!always14),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(sink_ready4),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~4 .extended_lut = "off";
defparam \sink_ready~4 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \sink_ready~4 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~5 (
	.dataa(!clr_break_line),
	.datab(!m0_write2),
	.datac(!mem_used_16),
	.datad(!wait_latency_counter_15),
	.datae(!wait_latency_counter_05),
	.dataf(!always15),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(sink_ready5),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~5 .extended_lut = "off";
defparam \sink_ready~5 .lut_mask = 64'hFFF7FFFDFFFFFFFF;
defparam \sink_ready~5 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~6 (
	.dataa(!clr_break_line),
	.datab(!m0_write2),
	.datac(!always16),
	.datad(!mem_used_17),
	.datae(!wait_latency_counter_16),
	.dataf(!wait_latency_counter_06),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(sink_ready6),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~6 .extended_lut = "off";
defparam \sink_ready~6 .lut_mask = 64'hFFFFFF7FFFFFFFDF;
defparam \sink_ready~6 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~7 (
	.dataa(!clr_break_line),
	.datab(!m0_write2),
	.datac(!mem_used_18),
	.datad(!wait_latency_counter_17),
	.datae(!wait_latency_counter_07),
	.dataf(!always17),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(sink_ready7),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~7 .extended_lut = "off";
defparam \sink_ready~7 .lut_mask = 64'hFFF7FFFDFFFFFFFF;
defparam \sink_ready~7 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~8 (
	.dataa(!clr_break_line),
	.datab(!m0_write2),
	.datac(!mem_used_19),
	.datad(!wait_latency_counter_18),
	.datae(!wait_latency_counter_08),
	.dataf(!always18),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(sink_ready8),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~8 .extended_lut = "off";
defparam \sink_ready~8 .lut_mask = 64'hFFF7FFFDFFFFFFFF;
defparam \sink_ready~8 .shared_arith = "off";

cyclonev_lcell_comb \WideOr0~6 (
	.dataa(!sink_ready),
	.datab(!sink_ready1),
	.datac(!sink_ready2),
	.datad(!\WideOr0~4_combout ),
	.datae(!\WideOr0~5_combout ),
	.dataf(!\sink_ready~9_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr01),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~6 .extended_lut = "off";
defparam \WideOr0~6 .lut_mask = 64'hFFFFFFFFFFFEFFFF;
defparam \WideOr0~6 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~10 (
	.dataa(!mem_used_14),
	.datab(!av_waitrequest_generated),
	.datac(!sink_ready3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(sink_ready9),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~10 .extended_lut = "off";
defparam \sink_ready~10 .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \sink_ready~10 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~11 (
	.dataa(!mem_used_15),
	.datab(!av_waitrequest_generated1),
	.datac(!sink_ready4),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(sink_ready10),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~11 .extended_lut = "off";
defparam \sink_ready~11 .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \sink_ready~11 .shared_arith = "off";

cyclonev_lcell_comb \src3_valid~0 (
	.dataa(!cp_valid),
	.datab(!src_channel_2),
	.datac(!src_channel_21),
	.datad(!Equal1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src3_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src3_valid~0 .extended_lut = "off";
defparam \src3_valid~0 .lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam \src3_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~12 (
	.dataa(!clr_break_line),
	.datab(!m0_write2),
	.datac(!mem_used_11),
	.datad(!wait_latency_counter_12),
	.datae(!wait_latency_counter_02),
	.dataf(!always11),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(sink_ready11),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~12 .extended_lut = "off";
defparam \sink_ready~12 .lut_mask = 64'hFFD7FF7DFFFFFFFF;
defparam \sink_ready~12 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~13 (
	.dataa(!clr_break_line),
	.datab(!m0_write2),
	.datac(!always12),
	.datad(!mem_used_12),
	.datae(!wait_latency_counter_13),
	.dataf(!wait_latency_counter_03),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(sink_ready12),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~13 .extended_lut = "off";
defparam \sink_ready~13 .lut_mask = 64'hFFFFDF7FFFFF7FDF;
defparam \sink_ready~13 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~14 (
	.dataa(!clr_break_line),
	.datab(!m0_write2),
	.datac(!always13),
	.datad(!mem_used_13),
	.datae(!wait_latency_counter_14),
	.dataf(!wait_latency_counter_04),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(sink_ready13),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~14 .extended_lut = "off";
defparam \sink_ready~14 .lut_mask = 64'hFFFFDF7FFFFF7FDF;
defparam \sink_ready~14 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~15 (
	.dataa(!clr_break_line),
	.datab(!m0_write2),
	.datac(!mem_used_16),
	.datad(!wait_latency_counter_15),
	.datae(!wait_latency_counter_05),
	.dataf(!always15),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(sink_ready14),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~15 .extended_lut = "off";
defparam \sink_ready~15 .lut_mask = 64'hFFD7FF7DFFFFFFFF;
defparam \sink_ready~15 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~16 (
	.dataa(!clr_break_line),
	.datab(!m0_write2),
	.datac(!always16),
	.datad(!mem_used_17),
	.datae(!wait_latency_counter_16),
	.dataf(!wait_latency_counter_06),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(sink_ready15),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~16 .extended_lut = "off";
defparam \sink_ready~16 .lut_mask = 64'hFFFFDF7FFFFF7FDF;
defparam \sink_ready~16 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~17 (
	.dataa(!clr_break_line),
	.datab(!m0_write2),
	.datac(!mem_used_18),
	.datad(!wait_latency_counter_17),
	.datae(!wait_latency_counter_07),
	.dataf(!always17),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(sink_ready16),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~17 .extended_lut = "off";
defparam \sink_ready~17 .lut_mask = 64'hFFD7FF7DFFFFFFFF;
defparam \sink_ready~17 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~18 (
	.dataa(!clr_break_line),
	.datab(!m0_write2),
	.datac(!mem_used_19),
	.datad(!wait_latency_counter_18),
	.datae(!wait_latency_counter_08),
	.dataf(!always18),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(sink_ready17),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~18 .extended_lut = "off";
defparam \sink_ready~18 .lut_mask = 64'hFFD7FF7DFFFFFFFF;
defparam \sink_ready~18 .shared_arith = "off";

cyclonev_lcell_comb \src2_valid~0 (
	.dataa(!cp_valid),
	.datab(!src_channel_2),
	.datac(!src_channel_21),
	.datad(!Equal1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src2_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src2_valid~0 .extended_lut = "off";
defparam \src2_valid~0 .lut_mask = 64'hF7FFF7FFF7FFF7FF;
defparam \src2_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \WideOr0~0 (
	.dataa(!wait_latency_counter_0),
	.datab(!wait_latency_counter_1),
	.datac(!m0_write),
	.datad(!m0_write2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~0 .extended_lut = "off";
defparam \WideOr0~0 .lut_mask = 64'hDFEFDFEFDFEFDFEF;
defparam \WideOr0~0 .shared_arith = "off";

cyclonev_lcell_comb \WideOr0~1 (
	.dataa(!mem_used_1),
	.datab(!saved_grant_0),
	.datac(!src_channel_2),
	.datad(!src_channel_21),
	.datae(!Equal1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~1 .extended_lut = "off";
defparam \WideOr0~1 .lut_mask = 64'hFFFFFFBFFFFFFFBF;
defparam \WideOr0~1 .shared_arith = "off";

cyclonev_lcell_comb \WideOr0~2 (
	.dataa(!wait_latency_counter_01),
	.datab(!wait_latency_counter_11),
	.datac(!m0_write1),
	.datad(!m0_write2),
	.datae(!write3),
	.dataf(!write4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~2 .extended_lut = "off";
defparam \WideOr0~2 .lut_mask = 64'hFFFFFFFFFFFFF7FB;
defparam \WideOr0~2 .shared_arith = "off";

cyclonev_lcell_comb \WideOr0~4 (
	.dataa(!mem_used_14),
	.datab(!av_waitrequest_generated),
	.datac(!sink_ready3),
	.datad(!mem_used_15),
	.datae(!av_waitrequest_generated1),
	.dataf(!sink_ready4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr0~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~4 .extended_lut = "off";
defparam \WideOr0~4 .lut_mask = 64'hFFBFFFFFFFFFFFFF;
defparam \WideOr0~4 .shared_arith = "off";

cyclonev_lcell_comb \WideOr0~5 (
	.dataa(!av_waitrequest),
	.datab(!av_waitrequest1),
	.datac(!sink_ready5),
	.datad(!sink_ready6),
	.datae(!sink_ready7),
	.dataf(!sink_ready8),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr0~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~5 .extended_lut = "off";
defparam \WideOr0~5 .lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam \WideOr0~5 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~9 (
	.dataa(!saved_grant_01),
	.datab(!write5),
	.datac(!src_channel_2),
	.datad(!src_channel_21),
	.datae(!Equal1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sink_ready~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~9 .extended_lut = "off";
defparam \sink_ready~9 .lut_mask = 64'hFF7FFFFFFF7FFFFF;
defparam \sink_ready~9 .shared_arith = "off";

endmodule

module first_nios2_system_first_nios2_system_mm_interconnect_0_cmd_demux_001 (
	clr_break_line,
	write,
	saved_grant_1,
	last_dest_id_2,
	has_pending_responses,
	i_read,
	Equal1,
	saved_grant_11,
	last_dest_id_3,
	read_latency_shift_reg,
	src1_valid,
	src0_valid,
	WideOr0)/* synthesis synthesis_greybox=1 */;
input 	clr_break_line;
input 	write;
input 	saved_grant_1;
input 	last_dest_id_2;
input 	has_pending_responses;
input 	i_read;
input 	Equal1;
input 	saved_grant_11;
input 	last_dest_id_3;
input 	read_latency_shift_reg;
output 	src1_valid;
output 	src0_valid;
output 	WideOr0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \src1_valid~0 (
	.dataa(!clr_break_line),
	.datab(!has_pending_responses),
	.datac(!i_read),
	.datad(!Equal1),
	.datae(!last_dest_id_3),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src1_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src1_valid~0 .extended_lut = "off";
defparam \src1_valid~0 .lut_mask = 64'hFFDFFFFFFFDFFFFF;
defparam \src1_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \src0_valid~0 (
	.dataa(!clr_break_line),
	.datab(!last_dest_id_2),
	.datac(!has_pending_responses),
	.datad(!i_read),
	.datae(!Equal1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src0_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src0_valid~0 .extended_lut = "off";
defparam \src0_valid~0 .lut_mask = 64'hF7FFFFFFF7FFFFFF;
defparam \src0_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \WideOr0~0 (
	.dataa(!write),
	.datab(!saved_grant_1),
	.datac(!Equal1),
	.datad(!saved_grant_11),
	.datae(!read_latency_shift_reg),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr0),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~0 .extended_lut = "off";
defparam \WideOr0~0 .lut_mask = 64'h53FFFFFF53FFFFFF;
defparam \WideOr0~0 .shared_arith = "off";

endmodule

module first_nios2_system_first_nios2_system_mm_interconnect_0_cmd_mux_002 (
	A_st_data_0,
	A_mem_baddr_4,
	A_mem_baddr_5,
	A_mem_baddr_8,
	A_mem_baddr_10,
	A_mem_baddr_9,
	A_mem_baddr_7,
	A_mem_baddr_6,
	clr_break_line,
	A_mem_baddr_3,
	A_mem_baddr_2,
	r_sync_rst,
	A_st_data_1,
	A_st_data_2,
	A_st_data_3,
	A_st_data_4,
	A_st_data_5,
	A_st_data_6,
	A_st_data_7,
	cp_valid,
	W_debug_mode,
	src_channel_2,
	src_channel_21,
	Equal1,
	saved_grant_0,
	write,
	saved_grant_1,
	last_dest_id_2,
	has_pending_responses,
	i_read,
	Equal11,
	WideOr11,
	src2_valid,
	src0_valid,
	src_payload,
	ic_fill_ap_offset_0,
	src_data_38,
	ic_fill_line_0,
	src_data_41,
	ic_fill_ap_offset_2,
	src_data_40,
	ic_fill_ap_offset_1,
	src_data_39,
	ic_fill_line_5,
	src_data_46,
	ic_fill_line_4,
	src_data_45,
	ic_fill_line_3,
	src_data_44,
	ic_fill_line_2,
	src_data_43,
	ic_fill_line_1,
	src_data_42,
	src_payload1,
	src_payload2,
	A_mem_byte_en_0,
	src_data_32,
	src_payload3,
	A_st_data_16,
	src_payload4,
	A_st_data_22,
	A_mem_byte_en_2,
	A_st_data_23,
	A_st_data_24,
	A_mem_byte_en_3,
	A_st_data_25,
	A_st_data_31,
	A_st_data_21,
	A_st_data_11,
	A_mem_byte_en_1,
	A_st_data_28,
	A_st_data_10,
	A_st_data_27,
	A_st_data_8,
	A_st_data_9,
	A_st_data_26,
	A_st_data_20,
	A_st_data_19,
	A_st_data_17,
	A_st_data_30,
	A_st_data_18,
	A_st_data_15,
	A_st_data_12,
	A_st_data_13,
	A_st_data_14,
	A_st_data_29,
	src_payload5,
	src_payload6,
	src_data_34,
	src_payload7,
	src_payload8,
	src_payload9,
	src_payload10,
	src_payload11,
	src_payload12,
	src_payload13,
	src_payload14,
	src_payload15,
	src_data_35,
	src_payload16,
	src_payload17,
	src_payload18,
	src_payload19,
	src_payload20,
	src_payload21,
	src_payload22,
	src_data_33,
	src_payload23,
	src_payload24,
	src_payload25,
	src_payload26,
	src_payload27,
	src_payload28,
	src_payload29,
	src_payload30,
	src_payload31,
	src_payload32,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	A_st_data_0;
input 	A_mem_baddr_4;
input 	A_mem_baddr_5;
input 	A_mem_baddr_8;
input 	A_mem_baddr_10;
input 	A_mem_baddr_9;
input 	A_mem_baddr_7;
input 	A_mem_baddr_6;
input 	clr_break_line;
input 	A_mem_baddr_3;
input 	A_mem_baddr_2;
input 	r_sync_rst;
input 	A_st_data_1;
input 	A_st_data_2;
input 	A_st_data_3;
input 	A_st_data_4;
input 	A_st_data_5;
input 	A_st_data_6;
input 	A_st_data_7;
input 	cp_valid;
input 	W_debug_mode;
input 	src_channel_2;
input 	src_channel_21;
input 	Equal1;
output 	saved_grant_0;
input 	write;
output 	saved_grant_1;
input 	last_dest_id_2;
input 	has_pending_responses;
input 	i_read;
input 	Equal11;
output 	WideOr11;
input 	src2_valid;
input 	src0_valid;
output 	src_payload;
input 	ic_fill_ap_offset_0;
output 	src_data_38;
input 	ic_fill_line_0;
output 	src_data_41;
input 	ic_fill_ap_offset_2;
output 	src_data_40;
input 	ic_fill_ap_offset_1;
output 	src_data_39;
input 	ic_fill_line_5;
output 	src_data_46;
input 	ic_fill_line_4;
output 	src_data_45;
input 	ic_fill_line_3;
output 	src_data_44;
input 	ic_fill_line_2;
output 	src_data_43;
input 	ic_fill_line_1;
output 	src_data_42;
output 	src_payload1;
output 	src_payload2;
input 	A_mem_byte_en_0;
output 	src_data_32;
output 	src_payload3;
input 	A_st_data_16;
output 	src_payload4;
input 	A_st_data_22;
input 	A_mem_byte_en_2;
input 	A_st_data_23;
input 	A_st_data_24;
input 	A_mem_byte_en_3;
input 	A_st_data_25;
input 	A_st_data_31;
input 	A_st_data_21;
input 	A_st_data_11;
input 	A_mem_byte_en_1;
input 	A_st_data_28;
input 	A_st_data_10;
input 	A_st_data_27;
input 	A_st_data_8;
input 	A_st_data_9;
input 	A_st_data_26;
input 	A_st_data_20;
input 	A_st_data_19;
input 	A_st_data_17;
input 	A_st_data_30;
input 	A_st_data_18;
input 	A_st_data_15;
input 	A_st_data_12;
input 	A_st_data_13;
input 	A_st_data_14;
input 	A_st_data_29;
output 	src_payload5;
output 	src_payload6;
output 	src_data_34;
output 	src_payload7;
output 	src_payload8;
output 	src_payload9;
output 	src_payload10;
output 	src_payload11;
output 	src_payload12;
output 	src_payload13;
output 	src_payload14;
output 	src_payload15;
output 	src_data_35;
output 	src_payload16;
output 	src_payload17;
output 	src_payload18;
output 	src_payload19;
output 	src_payload20;
output 	src_payload21;
output 	src_payload22;
output 	src_data_33;
output 	src_payload23;
output 	src_payload24;
output 	src_payload25;
output 	src_payload26;
output 	src_payload27;
output 	src_payload28;
output 	src_payload29;
output 	src_payload30;
output 	src_payload31;
output 	src_payload32;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \arb|grant[0]~0_combout ;
wire \arb|grant[1]~1_combout ;
wire \packet_in_progress~0_combout ;
wire \packet_in_progress~q ;
wire \update_grant~0_combout ;
wire \src_valid~0_combout ;


first_nios2_system_altera_merlin_arbitrator arb(
	.reset(r_sync_rst),
	.saved_grant_0(saved_grant_0),
	.write(write),
	.saved_grant_1(saved_grant_1),
	.src2_valid(src2_valid),
	.src0_valid(src0_valid),
	.grant_0(\arb|grant[0]~0_combout ),
	.packet_in_progress(\packet_in_progress~q ),
	.grant_1(\arb|grant[1]~1_combout ),
	.clk(clk_clk));

dffeas \saved_grant[0] (
	.clk(clk_clk),
	.d(\arb|grant[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~0_combout ),
	.q(saved_grant_0),
	.prn(vcc));
defparam \saved_grant[0] .is_wysiwyg = "true";
defparam \saved_grant[0] .power_up = "low";

dffeas \saved_grant[1] (
	.clk(clk_clk),
	.d(\arb|grant[1]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~0_combout ),
	.q(saved_grant_1),
	.prn(vcc));
defparam \saved_grant[1] .is_wysiwyg = "true";
defparam \saved_grant[1] .power_up = "low";

cyclonev_lcell_comb WideOr1(
	.dataa(!cp_valid),
	.datab(!saved_grant_0),
	.datac(!src_channel_2),
	.datad(!src_channel_21),
	.datae(!Equal1),
	.dataf(!\src_valid~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr11),
	.sumout(),
	.cout(),
	.shareout());
defparam WideOr1.extended_lut = "off";
defparam WideOr1.lut_mask = 64'hFFFFFFFFFFFFFEFF;
defparam WideOr1.shared_arith = "off";

cyclonev_lcell_comb \src_payload~0 (
	.dataa(!A_st_data_3),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~0 .extended_lut = "off";
defparam \src_payload~0 .lut_mask = 64'h7777777777777777;
defparam \src_payload~0 .shared_arith = "off";

cyclonev_lcell_comb \src_data[38] (
	.dataa(!A_mem_baddr_2),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!ic_fill_ap_offset_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_38),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[38] .extended_lut = "off";
defparam \src_data[38] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[38] .shared_arith = "off";

cyclonev_lcell_comb \src_data[41] (
	.dataa(!A_mem_baddr_5),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!ic_fill_line_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_41),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[41] .extended_lut = "off";
defparam \src_data[41] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[41] .shared_arith = "off";

cyclonev_lcell_comb \src_data[40] (
	.dataa(!A_mem_baddr_4),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!ic_fill_ap_offset_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_40),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[40] .extended_lut = "off";
defparam \src_data[40] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[40] .shared_arith = "off";

cyclonev_lcell_comb \src_data[39] (
	.dataa(!A_mem_baddr_3),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!ic_fill_ap_offset_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_39),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[39] .extended_lut = "off";
defparam \src_data[39] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[39] .shared_arith = "off";

cyclonev_lcell_comb \src_data[46] (
	.dataa(!A_mem_baddr_10),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!ic_fill_line_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_46),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[46] .extended_lut = "off";
defparam \src_data[46] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[46] .shared_arith = "off";

cyclonev_lcell_comb \src_data[45] (
	.dataa(!A_mem_baddr_9),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!ic_fill_line_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_45),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[45] .extended_lut = "off";
defparam \src_data[45] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[45] .shared_arith = "off";

cyclonev_lcell_comb \src_data[44] (
	.dataa(!A_mem_baddr_8),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!ic_fill_line_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_44),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[44] .extended_lut = "off";
defparam \src_data[44] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[44] .shared_arith = "off";

cyclonev_lcell_comb \src_data[43] (
	.dataa(!A_mem_baddr_7),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!ic_fill_line_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_43),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[43] .extended_lut = "off";
defparam \src_data[43] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[43] .shared_arith = "off";

cyclonev_lcell_comb \src_data[42] (
	.dataa(!A_mem_baddr_6),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!ic_fill_line_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_42),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[42] .extended_lut = "off";
defparam \src_data[42] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[42] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~1 (
	.dataa(!W_debug_mode),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~1 .extended_lut = "off";
defparam \src_payload~1 .lut_mask = 64'h7777777777777777;
defparam \src_payload~1 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~2 (
	.dataa(!A_st_data_0),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload2),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~2 .extended_lut = "off";
defparam \src_payload~2 .lut_mask = 64'h7777777777777777;
defparam \src_payload~2 .shared_arith = "off";

cyclonev_lcell_comb \src_data[32] (
	.dataa(!saved_grant_0),
	.datab(!saved_grant_1),
	.datac(!A_mem_byte_en_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_32),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[32] .extended_lut = "off";
defparam \src_data[32] .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \src_data[32] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~3 (
	.dataa(!A_st_data_1),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload3),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~3 .extended_lut = "off";
defparam \src_payload~3 .lut_mask = 64'h7777777777777777;
defparam \src_payload~3 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~4 (
	.dataa(!saved_grant_0),
	.datab(!A_st_data_16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload4),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~4 .extended_lut = "off";
defparam \src_payload~4 .lut_mask = 64'h7777777777777777;
defparam \src_payload~4 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~5 (
	.dataa(!A_st_data_2),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload5),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~5 .extended_lut = "off";
defparam \src_payload~5 .lut_mask = 64'h7777777777777777;
defparam \src_payload~5 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~6 (
	.dataa(!saved_grant_0),
	.datab(!A_st_data_20),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload6),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~6 .extended_lut = "off";
defparam \src_payload~6 .lut_mask = 64'h7777777777777777;
defparam \src_payload~6 .shared_arith = "off";

cyclonev_lcell_comb \src_data[34] (
	.dataa(!saved_grant_0),
	.datab(!saved_grant_1),
	.datac(!A_mem_byte_en_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_34),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[34] .extended_lut = "off";
defparam \src_data[34] .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \src_data[34] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~7 (
	.dataa(!saved_grant_0),
	.datab(!A_st_data_19),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload7),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~7 .extended_lut = "off";
defparam \src_payload~7 .lut_mask = 64'h7777777777777777;
defparam \src_payload~7 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~8 (
	.dataa(!saved_grant_0),
	.datab(!A_st_data_21),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload8),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~8 .extended_lut = "off";
defparam \src_payload~8 .lut_mask = 64'h7777777777777777;
defparam \src_payload~8 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~9 (
	.dataa(!saved_grant_0),
	.datab(!A_st_data_18),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload9),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~9 .extended_lut = "off";
defparam \src_payload~9 .lut_mask = 64'h7777777777777777;
defparam \src_payload~9 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~10 (
	.dataa(!saved_grant_0),
	.datab(!A_st_data_17),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload10),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~10 .extended_lut = "off";
defparam \src_payload~10 .lut_mask = 64'h7777777777777777;
defparam \src_payload~10 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~11 (
	.dataa(!A_st_data_4),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload11),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~11 .extended_lut = "off";
defparam \src_payload~11 .lut_mask = 64'h7777777777777777;
defparam \src_payload~11 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~12 (
	.dataa(!A_st_data_5),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload12),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~12 .extended_lut = "off";
defparam \src_payload~12 .lut_mask = 64'h7777777777777777;
defparam \src_payload~12 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~13 (
	.dataa(!A_st_data_6),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload13),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~13 .extended_lut = "off";
defparam \src_payload~13 .lut_mask = 64'h7777777777777777;
defparam \src_payload~13 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~14 (
	.dataa(!A_st_data_7),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload14),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~14 .extended_lut = "off";
defparam \src_payload~14 .lut_mask = 64'h7777777777777777;
defparam \src_payload~14 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~15 (
	.dataa(!saved_grant_0),
	.datab(!A_st_data_24),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload15),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~15 .extended_lut = "off";
defparam \src_payload~15 .lut_mask = 64'h7777777777777777;
defparam \src_payload~15 .shared_arith = "off";

cyclonev_lcell_comb \src_data[35] (
	.dataa(!saved_grant_0),
	.datab(!saved_grant_1),
	.datac(!A_mem_byte_en_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_35),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[35] .extended_lut = "off";
defparam \src_data[35] .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \src_data[35] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~16 (
	.dataa(!saved_grant_0),
	.datab(!A_st_data_25),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload16),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~16 .extended_lut = "off";
defparam \src_payload~16 .lut_mask = 64'h7777777777777777;
defparam \src_payload~16 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~17 (
	.dataa(!saved_grant_0),
	.datab(!A_st_data_26),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload17),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~17 .extended_lut = "off";
defparam \src_payload~17 .lut_mask = 64'h7777777777777777;
defparam \src_payload~17 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~18 (
	.dataa(!saved_grant_0),
	.datab(!A_st_data_27),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload18),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~18 .extended_lut = "off";
defparam \src_payload~18 .lut_mask = 64'h7777777777777777;
defparam \src_payload~18 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~19 (
	.dataa(!saved_grant_0),
	.datab(!A_st_data_22),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload19),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~19 .extended_lut = "off";
defparam \src_payload~19 .lut_mask = 64'h7777777777777777;
defparam \src_payload~19 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~20 (
	.dataa(!saved_grant_0),
	.datab(!A_st_data_23),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload20),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~20 .extended_lut = "off";
defparam \src_payload~20 .lut_mask = 64'h7777777777777777;
defparam \src_payload~20 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~21 (
	.dataa(!saved_grant_0),
	.datab(!A_st_data_31),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload21),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~21 .extended_lut = "off";
defparam \src_payload~21 .lut_mask = 64'h7777777777777777;
defparam \src_payload~21 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~22 (
	.dataa(!saved_grant_0),
	.datab(!A_st_data_11),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload22),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~22 .extended_lut = "off";
defparam \src_payload~22 .lut_mask = 64'h7777777777777777;
defparam \src_payload~22 .shared_arith = "off";

cyclonev_lcell_comb \src_data[33] (
	.dataa(!saved_grant_0),
	.datab(!saved_grant_1),
	.datac(!A_mem_byte_en_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_33),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[33] .extended_lut = "off";
defparam \src_data[33] .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \src_data[33] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~23 (
	.dataa(!saved_grant_0),
	.datab(!A_st_data_28),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload23),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~23 .extended_lut = "off";
defparam \src_payload~23 .lut_mask = 64'h7777777777777777;
defparam \src_payload~23 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~24 (
	.dataa(!saved_grant_0),
	.datab(!A_st_data_10),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload24),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~24 .extended_lut = "off";
defparam \src_payload~24 .lut_mask = 64'h7777777777777777;
defparam \src_payload~24 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~25 (
	.dataa(!saved_grant_0),
	.datab(!A_st_data_8),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload25),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~25 .extended_lut = "off";
defparam \src_payload~25 .lut_mask = 64'h7777777777777777;
defparam \src_payload~25 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~26 (
	.dataa(!saved_grant_0),
	.datab(!A_st_data_9),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload26),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~26 .extended_lut = "off";
defparam \src_payload~26 .lut_mask = 64'h7777777777777777;
defparam \src_payload~26 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~27 (
	.dataa(!saved_grant_0),
	.datab(!A_st_data_30),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload27),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~27 .extended_lut = "off";
defparam \src_payload~27 .lut_mask = 64'h7777777777777777;
defparam \src_payload~27 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~28 (
	.dataa(!saved_grant_0),
	.datab(!A_st_data_15),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload28),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~28 .extended_lut = "off";
defparam \src_payload~28 .lut_mask = 64'h7777777777777777;
defparam \src_payload~28 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~29 (
	.dataa(!saved_grant_0),
	.datab(!A_st_data_12),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload29),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~29 .extended_lut = "off";
defparam \src_payload~29 .lut_mask = 64'h7777777777777777;
defparam \src_payload~29 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~30 (
	.dataa(!saved_grant_0),
	.datab(!A_st_data_13),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload30),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~30 .extended_lut = "off";
defparam \src_payload~30 .lut_mask = 64'h7777777777777777;
defparam \src_payload~30 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~31 (
	.dataa(!saved_grant_0),
	.datab(!A_st_data_14),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload31),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~31 .extended_lut = "off";
defparam \src_payload~31 .lut_mask = 64'h7777777777777777;
defparam \src_payload~31 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~32 (
	.dataa(!saved_grant_0),
	.datab(!A_st_data_29),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload32),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~32 .extended_lut = "off";
defparam \src_payload~32 .lut_mask = 64'h7777777777777777;
defparam \src_payload~32 .shared_arith = "off";

cyclonev_lcell_comb \packet_in_progress~0 (
	.dataa(!\update_grant~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\packet_in_progress~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \packet_in_progress~0 .extended_lut = "off";
defparam \packet_in_progress~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \packet_in_progress~0 .shared_arith = "off";

dffeas packet_in_progress(
	.clk(clk_clk),
	.d(\packet_in_progress~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\packet_in_progress~q ),
	.prn(vcc));
defparam packet_in_progress.is_wysiwyg = "true";
defparam packet_in_progress.power_up = "low";

cyclonev_lcell_comb \update_grant~0 (
	.dataa(!saved_grant_0),
	.datab(!write),
	.datac(!saved_grant_1),
	.datad(!WideOr11),
	.datae(!\packet_in_progress~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\update_grant~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \update_grant~0 .extended_lut = "off";
defparam \update_grant~0 .lut_mask = 64'hFF7F3F7FFF7F3F7F;
defparam \update_grant~0 .shared_arith = "off";

cyclonev_lcell_comb \src_valid~0 (
	.dataa(!clr_break_line),
	.datab(!saved_grant_1),
	.datac(!last_dest_id_2),
	.datad(!has_pending_responses),
	.datae(!i_read),
	.dataf(!Equal11),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_valid~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_valid~0 .extended_lut = "off";
defparam \src_valid~0 .lut_mask = 64'hFF7FFFFFFFFFFFFF;
defparam \src_valid~0 .shared_arith = "off";

endmodule

module first_nios2_system_altera_merlin_arbitrator (
	reset,
	saved_grant_0,
	write,
	saved_grant_1,
	src2_valid,
	src0_valid,
	grant_0,
	packet_in_progress,
	grant_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	saved_grant_0;
input 	write;
input 	saved_grant_1;
input 	src2_valid;
input 	src0_valid;
output 	grant_0;
input 	packet_in_progress;
output 	grant_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \top_priority_reg[0]~1_combout ;
wire \top_priority_reg[0]~0_combout ;
wire \top_priority_reg[0]~q ;
wire \top_priority_reg[1]~q ;


cyclonev_lcell_comb \grant[0]~0 (
	.dataa(!src2_valid),
	.datab(!src0_valid),
	.datac(!\top_priority_reg[0]~q ),
	.datad(!\top_priority_reg[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(grant_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \grant[0]~0 .extended_lut = "off";
defparam \grant[0]~0 .lut_mask = 64'hFDFFFDFFFDFFFDFF;
defparam \grant[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \grant[1]~1 (
	.dataa(!src2_valid),
	.datab(!src0_valid),
	.datac(!\top_priority_reg[0]~q ),
	.datad(!\top_priority_reg[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(grant_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \grant[1]~1 .extended_lut = "off";
defparam \grant[1]~1 .lut_mask = 64'hFBFFFBFFFBFFFBFF;
defparam \grant[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \top_priority_reg[0]~1 (
	.dataa(!grant_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~1 .extended_lut = "off";
defparam \top_priority_reg[0]~1 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \top_priority_reg[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \top_priority_reg[0]~0 (
	.dataa(!saved_grant_0),
	.datab(!write),
	.datac(!src2_valid),
	.datad(!saved_grant_1),
	.datae(!src0_valid),
	.dataf(!packet_in_progress),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~0 .extended_lut = "off";
defparam \top_priority_reg[0]~0 .lut_mask = 64'hFFFFFFFF7BB7B77B;
defparam \top_priority_reg[0]~0 .shared_arith = "off";

dffeas \top_priority_reg[0] (
	.clk(clk),
	.d(\top_priority_reg[0]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~0_combout ),
	.q(\top_priority_reg[0]~q ),
	.prn(vcc));
defparam \top_priority_reg[0] .is_wysiwyg = "true";
defparam \top_priority_reg[0] .power_up = "low";

dffeas \top_priority_reg[1] (
	.clk(clk),
	.d(grant_0),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~0_combout ),
	.q(\top_priority_reg[1]~q ),
	.prn(vcc));
defparam \top_priority_reg[1] .is_wysiwyg = "true";
defparam \top_priority_reg[1] .power_up = "low";

endmodule

module first_nios2_system_first_nios2_system_mm_interconnect_0_cmd_mux_002_1 (
	A_st_data_0,
	A_mem_baddr_4,
	A_mem_baddr_5,
	A_mem_baddr_8,
	A_mem_baddr_14,
	A_mem_baddr_13,
	A_mem_baddr_12,
	A_mem_baddr_11,
	A_mem_baddr_10,
	A_mem_baddr_9,
	A_mem_baddr_7,
	A_mem_baddr_6,
	clr_break_line,
	A_mem_baddr_3,
	A_mem_baddr_2,
	r_sync_rst,
	A_st_data_1,
	A_st_data_2,
	A_st_data_3,
	A_st_data_4,
	A_st_data_5,
	A_st_data_6,
	A_st_data_7,
	cp_valid,
	saved_grant_0,
	src_channel_2,
	src_channel_21,
	Equal1,
	has_pending_responses,
	i_read,
	ic_fill_tag_3,
	ic_fill_tag_2,
	ic_fill_tag_1,
	ic_fill_tag_0,
	Equal11,
	saved_grant_1,
	last_dest_id_3,
	WideOr11,
	read_latency_shift_reg,
	src3_valid,
	src1_valid,
	ic_fill_ap_offset_0,
	ic_fill_line_0,
	ic_fill_ap_offset_2,
	ic_fill_ap_offset_1,
	ic_fill_line_5,
	ic_fill_line_4,
	ic_fill_line_3,
	ic_fill_line_2,
	ic_fill_line_1,
	A_mem_byte_en_0,
	src_payload,
	src_data_38,
	src_data_39,
	src_data_40,
	src_data_41,
	src_data_42,
	src_data_43,
	src_data_44,
	src_data_45,
	src_data_46,
	src_data_47,
	src_data_48,
	src_data_49,
	src_data_50,
	src_data_32,
	A_st_data_16,
	src_payload1,
	src_payload2,
	src_payload3,
	src_payload4,
	src_payload5,
	src_payload6,
	src_payload7,
	A_st_data_22,
	src_payload8,
	A_mem_byte_en_2,
	src_data_34,
	A_st_data_23,
	src_payload9,
	A_st_data_24,
	src_payload10,
	A_mem_byte_en_3,
	src_data_35,
	A_st_data_25,
	src_payload11,
	A_st_data_31,
	src_payload12,
	A_st_data_21,
	src_payload13,
	A_st_data_11,
	src_payload14,
	A_mem_byte_en_1,
	src_data_33,
	A_st_data_28,
	src_payload15,
	A_st_data_10,
	src_payload16,
	A_st_data_27,
	src_payload17,
	A_st_data_8,
	src_payload18,
	A_st_data_9,
	src_payload19,
	A_st_data_26,
	src_payload20,
	A_st_data_20,
	src_payload21,
	A_st_data_19,
	src_payload22,
	A_st_data_17,
	src_payload23,
	A_st_data_30,
	src_payload24,
	A_st_data_18,
	src_payload25,
	src_payload26,
	A_st_data_15,
	src_payload27,
	A_st_data_12,
	src_payload28,
	A_st_data_13,
	src_payload29,
	A_st_data_14,
	src_payload30,
	A_st_data_29,
	src_payload31,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	A_st_data_0;
input 	A_mem_baddr_4;
input 	A_mem_baddr_5;
input 	A_mem_baddr_8;
input 	A_mem_baddr_14;
input 	A_mem_baddr_13;
input 	A_mem_baddr_12;
input 	A_mem_baddr_11;
input 	A_mem_baddr_10;
input 	A_mem_baddr_9;
input 	A_mem_baddr_7;
input 	A_mem_baddr_6;
input 	clr_break_line;
input 	A_mem_baddr_3;
input 	A_mem_baddr_2;
input 	r_sync_rst;
input 	A_st_data_1;
input 	A_st_data_2;
input 	A_st_data_3;
input 	A_st_data_4;
input 	A_st_data_5;
input 	A_st_data_6;
input 	A_st_data_7;
input 	cp_valid;
output 	saved_grant_0;
input 	src_channel_2;
input 	src_channel_21;
input 	Equal1;
input 	has_pending_responses;
input 	i_read;
input 	ic_fill_tag_3;
input 	ic_fill_tag_2;
input 	ic_fill_tag_1;
input 	ic_fill_tag_0;
input 	Equal11;
output 	saved_grant_1;
input 	last_dest_id_3;
output 	WideOr11;
input 	read_latency_shift_reg;
input 	src3_valid;
input 	src1_valid;
input 	ic_fill_ap_offset_0;
input 	ic_fill_line_0;
input 	ic_fill_ap_offset_2;
input 	ic_fill_ap_offset_1;
input 	ic_fill_line_5;
input 	ic_fill_line_4;
input 	ic_fill_line_3;
input 	ic_fill_line_2;
input 	ic_fill_line_1;
input 	A_mem_byte_en_0;
output 	src_payload;
output 	src_data_38;
output 	src_data_39;
output 	src_data_40;
output 	src_data_41;
output 	src_data_42;
output 	src_data_43;
output 	src_data_44;
output 	src_data_45;
output 	src_data_46;
output 	src_data_47;
output 	src_data_48;
output 	src_data_49;
output 	src_data_50;
output 	src_data_32;
input 	A_st_data_16;
output 	src_payload1;
output 	src_payload2;
output 	src_payload3;
output 	src_payload4;
output 	src_payload5;
output 	src_payload6;
output 	src_payload7;
input 	A_st_data_22;
output 	src_payload8;
input 	A_mem_byte_en_2;
output 	src_data_34;
input 	A_st_data_23;
output 	src_payload9;
input 	A_st_data_24;
output 	src_payload10;
input 	A_mem_byte_en_3;
output 	src_data_35;
input 	A_st_data_25;
output 	src_payload11;
input 	A_st_data_31;
output 	src_payload12;
input 	A_st_data_21;
output 	src_payload13;
input 	A_st_data_11;
output 	src_payload14;
input 	A_mem_byte_en_1;
output 	src_data_33;
input 	A_st_data_28;
output 	src_payload15;
input 	A_st_data_10;
output 	src_payload16;
input 	A_st_data_27;
output 	src_payload17;
input 	A_st_data_8;
output 	src_payload18;
input 	A_st_data_9;
output 	src_payload19;
input 	A_st_data_26;
output 	src_payload20;
input 	A_st_data_20;
output 	src_payload21;
input 	A_st_data_19;
output 	src_payload22;
input 	A_st_data_17;
output 	src_payload23;
input 	A_st_data_30;
output 	src_payload24;
input 	A_st_data_18;
output 	src_payload25;
output 	src_payload26;
input 	A_st_data_15;
output 	src_payload27;
input 	A_st_data_12;
output 	src_payload28;
input 	A_st_data_13;
output 	src_payload29;
input 	A_st_data_14;
output 	src_payload30;
input 	A_st_data_29;
output 	src_payload31;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \arb|grant[0]~0_combout ;
wire \arb|grant[1]~1_combout ;
wire \packet_in_progress~0_combout ;
wire \packet_in_progress~q ;
wire \update_grant~0_combout ;
wire \src_valid~0_combout ;


first_nios2_system_altera_merlin_arbitrator_1 arb(
	.reset(r_sync_rst),
	.saved_grant_0(saved_grant_0),
	.saved_grant_1(saved_grant_1),
	.read_latency_shift_reg(read_latency_shift_reg),
	.src3_valid(src3_valid),
	.src1_valid(src1_valid),
	.grant_0(\arb|grant[0]~0_combout ),
	.packet_in_progress(\packet_in_progress~q ),
	.grant_1(\arb|grant[1]~1_combout ),
	.clk(clk_clk));

dffeas \saved_grant[0] (
	.clk(clk_clk),
	.d(\arb|grant[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~0_combout ),
	.q(saved_grant_0),
	.prn(vcc));
defparam \saved_grant[0] .is_wysiwyg = "true";
defparam \saved_grant[0] .power_up = "low";

dffeas \saved_grant[1] (
	.clk(clk_clk),
	.d(\arb|grant[1]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~0_combout ),
	.q(saved_grant_1),
	.prn(vcc));
defparam \saved_grant[1] .is_wysiwyg = "true";
defparam \saved_grant[1] .power_up = "low";

cyclonev_lcell_comb WideOr1(
	.dataa(!cp_valid),
	.datab(!saved_grant_0),
	.datac(!src_channel_2),
	.datad(!src_channel_21),
	.datae(!Equal1),
	.dataf(!\src_valid~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr11),
	.sumout(),
	.cout(),
	.shareout());
defparam WideOr1.extended_lut = "off";
defparam WideOr1.lut_mask = 64'hFFFFFFFFFEFFFFFF;
defparam WideOr1.shared_arith = "off";

cyclonev_lcell_comb \src_payload~0 (
	.dataa(!A_st_data_0),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~0 .extended_lut = "off";
defparam \src_payload~0 .lut_mask = 64'h7777777777777777;
defparam \src_payload~0 .shared_arith = "off";

cyclonev_lcell_comb \src_data[38] (
	.dataa(!A_mem_baddr_2),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!ic_fill_ap_offset_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_38),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[38] .extended_lut = "off";
defparam \src_data[38] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[38] .shared_arith = "off";

cyclonev_lcell_comb \src_data[39] (
	.dataa(!A_mem_baddr_3),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!ic_fill_ap_offset_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_39),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[39] .extended_lut = "off";
defparam \src_data[39] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[39] .shared_arith = "off";

cyclonev_lcell_comb \src_data[40] (
	.dataa(!A_mem_baddr_4),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!ic_fill_ap_offset_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_40),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[40] .extended_lut = "off";
defparam \src_data[40] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[40] .shared_arith = "off";

cyclonev_lcell_comb \src_data[41] (
	.dataa(!A_mem_baddr_5),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!ic_fill_line_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_41),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[41] .extended_lut = "off";
defparam \src_data[41] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[41] .shared_arith = "off";

cyclonev_lcell_comb \src_data[42] (
	.dataa(!A_mem_baddr_6),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!ic_fill_line_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_42),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[42] .extended_lut = "off";
defparam \src_data[42] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[42] .shared_arith = "off";

cyclonev_lcell_comb \src_data[43] (
	.dataa(!A_mem_baddr_7),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!ic_fill_line_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_43),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[43] .extended_lut = "off";
defparam \src_data[43] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[43] .shared_arith = "off";

cyclonev_lcell_comb \src_data[44] (
	.dataa(!A_mem_baddr_8),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!ic_fill_line_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_44),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[44] .extended_lut = "off";
defparam \src_data[44] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[44] .shared_arith = "off";

cyclonev_lcell_comb \src_data[45] (
	.dataa(!A_mem_baddr_9),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!ic_fill_line_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_45),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[45] .extended_lut = "off";
defparam \src_data[45] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[45] .shared_arith = "off";

cyclonev_lcell_comb \src_data[46] (
	.dataa(!A_mem_baddr_10),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!ic_fill_line_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_46),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[46] .extended_lut = "off";
defparam \src_data[46] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[46] .shared_arith = "off";

cyclonev_lcell_comb \src_data[47] (
	.dataa(!A_mem_baddr_11),
	.datab(!saved_grant_0),
	.datac(!ic_fill_tag_0),
	.datad(!saved_grant_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_47),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[47] .extended_lut = "off";
defparam \src_data[47] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[47] .shared_arith = "off";

cyclonev_lcell_comb \src_data[48] (
	.dataa(!A_mem_baddr_12),
	.datab(!saved_grant_0),
	.datac(!ic_fill_tag_1),
	.datad(!saved_grant_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_48),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[48] .extended_lut = "off";
defparam \src_data[48] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[48] .shared_arith = "off";

cyclonev_lcell_comb \src_data[49] (
	.dataa(!A_mem_baddr_13),
	.datab(!saved_grant_0),
	.datac(!ic_fill_tag_2),
	.datad(!saved_grant_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_49),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[49] .extended_lut = "off";
defparam \src_data[49] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[49] .shared_arith = "off";

cyclonev_lcell_comb \src_data[50] (
	.dataa(!A_mem_baddr_14),
	.datab(!saved_grant_0),
	.datac(!ic_fill_tag_3),
	.datad(!saved_grant_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_50),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[50] .extended_lut = "off";
defparam \src_data[50] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[50] .shared_arith = "off";

cyclonev_lcell_comb \src_data[32] (
	.dataa(!saved_grant_0),
	.datab(!saved_grant_1),
	.datac(!A_mem_byte_en_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_32),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[32] .extended_lut = "off";
defparam \src_data[32] .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \src_data[32] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~1 (
	.dataa(!A_st_data_1),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~1 .extended_lut = "off";
defparam \src_payload~1 .lut_mask = 64'h7777777777777777;
defparam \src_payload~1 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~2 (
	.dataa(!A_st_data_2),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload2),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~2 .extended_lut = "off";
defparam \src_payload~2 .lut_mask = 64'h7777777777777777;
defparam \src_payload~2 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~3 (
	.dataa(!A_st_data_3),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload3),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~3 .extended_lut = "off";
defparam \src_payload~3 .lut_mask = 64'h7777777777777777;
defparam \src_payload~3 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~4 (
	.dataa(!A_st_data_4),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload4),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~4 .extended_lut = "off";
defparam \src_payload~4 .lut_mask = 64'h7777777777777777;
defparam \src_payload~4 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~5 (
	.dataa(!A_st_data_5),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload5),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~5 .extended_lut = "off";
defparam \src_payload~5 .lut_mask = 64'h7777777777777777;
defparam \src_payload~5 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~6 (
	.dataa(!A_st_data_6),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload6),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~6 .extended_lut = "off";
defparam \src_payload~6 .lut_mask = 64'h7777777777777777;
defparam \src_payload~6 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~7 (
	.dataa(!A_st_data_7),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload7),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~7 .extended_lut = "off";
defparam \src_payload~7 .lut_mask = 64'h7777777777777777;
defparam \src_payload~7 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~8 (
	.dataa(!saved_grant_0),
	.datab(!A_st_data_22),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload8),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~8 .extended_lut = "off";
defparam \src_payload~8 .lut_mask = 64'h7777777777777777;
defparam \src_payload~8 .shared_arith = "off";

cyclonev_lcell_comb \src_data[34] (
	.dataa(!saved_grant_0),
	.datab(!saved_grant_1),
	.datac(!A_mem_byte_en_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_34),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[34] .extended_lut = "off";
defparam \src_data[34] .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \src_data[34] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~9 (
	.dataa(!saved_grant_0),
	.datab(!A_st_data_23),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload9),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~9 .extended_lut = "off";
defparam \src_payload~9 .lut_mask = 64'h7777777777777777;
defparam \src_payload~9 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~10 (
	.dataa(!saved_grant_0),
	.datab(!A_st_data_24),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload10),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~10 .extended_lut = "off";
defparam \src_payload~10 .lut_mask = 64'h7777777777777777;
defparam \src_payload~10 .shared_arith = "off";

cyclonev_lcell_comb \src_data[35] (
	.dataa(!saved_grant_0),
	.datab(!saved_grant_1),
	.datac(!A_mem_byte_en_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_35),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[35] .extended_lut = "off";
defparam \src_data[35] .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \src_data[35] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~11 (
	.dataa(!saved_grant_0),
	.datab(!A_st_data_25),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload11),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~11 .extended_lut = "off";
defparam \src_payload~11 .lut_mask = 64'h7777777777777777;
defparam \src_payload~11 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~12 (
	.dataa(!saved_grant_0),
	.datab(!A_st_data_31),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload12),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~12 .extended_lut = "off";
defparam \src_payload~12 .lut_mask = 64'h7777777777777777;
defparam \src_payload~12 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~13 (
	.dataa(!saved_grant_0),
	.datab(!A_st_data_21),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload13),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~13 .extended_lut = "off";
defparam \src_payload~13 .lut_mask = 64'h7777777777777777;
defparam \src_payload~13 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~14 (
	.dataa(!saved_grant_0),
	.datab(!A_st_data_11),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload14),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~14 .extended_lut = "off";
defparam \src_payload~14 .lut_mask = 64'h7777777777777777;
defparam \src_payload~14 .shared_arith = "off";

cyclonev_lcell_comb \src_data[33] (
	.dataa(!saved_grant_0),
	.datab(!saved_grant_1),
	.datac(!A_mem_byte_en_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_33),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[33] .extended_lut = "off";
defparam \src_data[33] .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \src_data[33] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~15 (
	.dataa(!saved_grant_0),
	.datab(!A_st_data_28),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload15),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~15 .extended_lut = "off";
defparam \src_payload~15 .lut_mask = 64'h7777777777777777;
defparam \src_payload~15 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~16 (
	.dataa(!saved_grant_0),
	.datab(!A_st_data_10),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload16),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~16 .extended_lut = "off";
defparam \src_payload~16 .lut_mask = 64'h7777777777777777;
defparam \src_payload~16 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~17 (
	.dataa(!saved_grant_0),
	.datab(!A_st_data_27),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload17),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~17 .extended_lut = "off";
defparam \src_payload~17 .lut_mask = 64'h7777777777777777;
defparam \src_payload~17 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~18 (
	.dataa(!saved_grant_0),
	.datab(!A_st_data_8),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload18),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~18 .extended_lut = "off";
defparam \src_payload~18 .lut_mask = 64'h7777777777777777;
defparam \src_payload~18 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~19 (
	.dataa(!saved_grant_0),
	.datab(!A_st_data_9),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload19),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~19 .extended_lut = "off";
defparam \src_payload~19 .lut_mask = 64'h7777777777777777;
defparam \src_payload~19 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~20 (
	.dataa(!saved_grant_0),
	.datab(!A_st_data_26),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload20),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~20 .extended_lut = "off";
defparam \src_payload~20 .lut_mask = 64'h7777777777777777;
defparam \src_payload~20 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~21 (
	.dataa(!saved_grant_0),
	.datab(!A_st_data_20),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload21),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~21 .extended_lut = "off";
defparam \src_payload~21 .lut_mask = 64'h7777777777777777;
defparam \src_payload~21 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~22 (
	.dataa(!saved_grant_0),
	.datab(!A_st_data_19),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload22),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~22 .extended_lut = "off";
defparam \src_payload~22 .lut_mask = 64'h7777777777777777;
defparam \src_payload~22 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~23 (
	.dataa(!saved_grant_0),
	.datab(!A_st_data_17),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload23),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~23 .extended_lut = "off";
defparam \src_payload~23 .lut_mask = 64'h7777777777777777;
defparam \src_payload~23 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~24 (
	.dataa(!saved_grant_0),
	.datab(!A_st_data_30),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload24),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~24 .extended_lut = "off";
defparam \src_payload~24 .lut_mask = 64'h7777777777777777;
defparam \src_payload~24 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~25 (
	.dataa(!saved_grant_0),
	.datab(!A_st_data_18),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload25),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~25 .extended_lut = "off";
defparam \src_payload~25 .lut_mask = 64'h7777777777777777;
defparam \src_payload~25 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~26 (
	.dataa(!saved_grant_0),
	.datab(!A_st_data_16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload26),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~26 .extended_lut = "off";
defparam \src_payload~26 .lut_mask = 64'h7777777777777777;
defparam \src_payload~26 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~27 (
	.dataa(!saved_grant_0),
	.datab(!A_st_data_15),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload27),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~27 .extended_lut = "off";
defparam \src_payload~27 .lut_mask = 64'h7777777777777777;
defparam \src_payload~27 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~28 (
	.dataa(!saved_grant_0),
	.datab(!A_st_data_12),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload28),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~28 .extended_lut = "off";
defparam \src_payload~28 .lut_mask = 64'h7777777777777777;
defparam \src_payload~28 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~29 (
	.dataa(!saved_grant_0),
	.datab(!A_st_data_13),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload29),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~29 .extended_lut = "off";
defparam \src_payload~29 .lut_mask = 64'h7777777777777777;
defparam \src_payload~29 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~30 (
	.dataa(!saved_grant_0),
	.datab(!A_st_data_14),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload30),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~30 .extended_lut = "off";
defparam \src_payload~30 .lut_mask = 64'h7777777777777777;
defparam \src_payload~30 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~31 (
	.dataa(!saved_grant_0),
	.datab(!A_st_data_29),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload31),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~31 .extended_lut = "off";
defparam \src_payload~31 .lut_mask = 64'h7777777777777777;
defparam \src_payload~31 .shared_arith = "off";

cyclonev_lcell_comb \packet_in_progress~0 (
	.dataa(!\update_grant~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\packet_in_progress~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \packet_in_progress~0 .extended_lut = "off";
defparam \packet_in_progress~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \packet_in_progress~0 .shared_arith = "off";

dffeas packet_in_progress(
	.clk(clk_clk),
	.d(\packet_in_progress~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\packet_in_progress~q ),
	.prn(vcc));
defparam packet_in_progress.is_wysiwyg = "true";
defparam packet_in_progress.power_up = "low";

cyclonev_lcell_comb \update_grant~0 (
	.dataa(!saved_grant_0),
	.datab(!saved_grant_1),
	.datac(!WideOr11),
	.datad(!read_latency_shift_reg),
	.datae(!\packet_in_progress~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\update_grant~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \update_grant~0 .extended_lut = "off";
defparam \update_grant~0 .lut_mask = 64'hF7FF37FFF7FF37FF;
defparam \update_grant~0 .shared_arith = "off";

cyclonev_lcell_comb \src_valid~0 (
	.dataa(!clr_break_line),
	.datab(!has_pending_responses),
	.datac(!i_read),
	.datad(!Equal11),
	.datae(!saved_grant_1),
	.dataf(!last_dest_id_3),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_valid~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_valid~0 .extended_lut = "off";
defparam \src_valid~0 .lut_mask = 64'hFFDFFFFFFFFFFFFF;
defparam \src_valid~0 .shared_arith = "off";

endmodule

module first_nios2_system_altera_merlin_arbitrator_1 (
	reset,
	saved_grant_0,
	saved_grant_1,
	read_latency_shift_reg,
	src3_valid,
	src1_valid,
	grant_0,
	packet_in_progress,
	grant_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	saved_grant_0;
input 	saved_grant_1;
input 	read_latency_shift_reg;
input 	src3_valid;
input 	src1_valid;
output 	grant_0;
input 	packet_in_progress;
output 	grant_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \top_priority_reg[0]~1_combout ;
wire \top_priority_reg[0]~0_combout ;
wire \top_priority_reg[0]~q ;
wire \top_priority_reg[1]~q ;


cyclonev_lcell_comb \grant[0]~0 (
	.dataa(!src3_valid),
	.datab(!src1_valid),
	.datac(!\top_priority_reg[0]~q ),
	.datad(!\top_priority_reg[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(grant_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \grant[0]~0 .extended_lut = "off";
defparam \grant[0]~0 .lut_mask = 64'hFDFFFDFFFDFFFDFF;
defparam \grant[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \grant[1]~1 (
	.dataa(!src3_valid),
	.datab(!src1_valid),
	.datac(!\top_priority_reg[0]~q ),
	.datad(!\top_priority_reg[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(grant_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \grant[1]~1 .extended_lut = "off";
defparam \grant[1]~1 .lut_mask = 64'hFBFFFBFFFBFFFBFF;
defparam \grant[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \top_priority_reg[0]~1 (
	.dataa(!grant_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~1 .extended_lut = "off";
defparam \top_priority_reg[0]~1 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \top_priority_reg[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \top_priority_reg[0]~0 (
	.dataa(!saved_grant_0),
	.datab(!src3_valid),
	.datac(!saved_grant_1),
	.datad(!src1_valid),
	.datae(!read_latency_shift_reg),
	.dataf(!packet_in_progress),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~0 .extended_lut = "off";
defparam \top_priority_reg[0]~0 .lut_mask = 64'hFFFFFFFF6996FFFF;
defparam \top_priority_reg[0]~0 .shared_arith = "off";

dffeas \top_priority_reg[0] (
	.clk(clk),
	.d(\top_priority_reg[0]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~0_combout ),
	.q(\top_priority_reg[0]~q ),
	.prn(vcc));
defparam \top_priority_reg[0] .is_wysiwyg = "true";
defparam \top_priority_reg[0] .power_up = "low";

dffeas \top_priority_reg[1] (
	.clk(clk),
	.d(grant_0),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~0_combout ),
	.q(\top_priority_reg[1]~q ),
	.prn(vcc));
defparam \top_priority_reg[1] .is_wysiwyg = "true";
defparam \top_priority_reg[1] .power_up = "low";

endmodule

module first_nios2_system_first_nios2_system_mm_interconnect_0_router (
	A_mem_baddr_4,
	A_mem_baddr_5,
	A_mem_baddr_8,
	A_mem_baddr_16,
	A_mem_baddr_15,
	A_mem_baddr_14,
	A_mem_baddr_13,
	Equal1,
	A_mem_baddr_12,
	A_mem_baddr_11,
	A_mem_baddr_10,
	A_mem_baddr_9,
	Equal2,
	A_mem_baddr_7,
	A_mem_baddr_6,
	Equal15,
	A_mem_baddr_3,
	Equal14,
	Equal6,
	Equal61,
	always1,
	Equal16,
	Equal21,
	uav_read,
	Equal22,
	always11,
	always12,
	src_channel_2,
	src_channel_21,
	Equal11,
	always13,
	always14,
	always15,
	always16,
	always17,
	always18,
	always19,
	always110,
	always111)/* synthesis synthesis_greybox=1 */;
input 	A_mem_baddr_4;
input 	A_mem_baddr_5;
input 	A_mem_baddr_8;
input 	A_mem_baddr_16;
input 	A_mem_baddr_15;
input 	A_mem_baddr_14;
input 	A_mem_baddr_13;
output 	Equal1;
input 	A_mem_baddr_12;
input 	A_mem_baddr_11;
input 	A_mem_baddr_10;
input 	A_mem_baddr_9;
output 	Equal2;
input 	A_mem_baddr_7;
input 	A_mem_baddr_6;
output 	Equal15;
input 	A_mem_baddr_3;
output 	Equal14;
output 	Equal6;
output 	Equal61;
output 	always1;
output 	Equal16;
output 	Equal21;
input 	uav_read;
output 	Equal22;
output 	always11;
output 	always12;
output 	src_channel_2;
output 	src_channel_21;
output 	Equal11;
output 	always13;
output 	always14;
output 	always15;
output 	always16;
output 	always17;
output 	always18;
output 	always19;
output 	always110;
output 	always111;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Equal15~0_combout ;
wire \Equal15~2_combout ;
wire \src_channel[2]~0_combout ;
wire \src_channel[2]~1_combout ;
wire \Equal2~3_combout ;
wire \always1~8_combout ;
wire \always1~10_combout ;


cyclonev_lcell_comb \Equal1~0 (
	.dataa(!A_mem_baddr_16),
	.datab(!A_mem_baddr_15),
	.datac(!A_mem_baddr_14),
	.datad(!A_mem_baddr_13),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal1),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal1~0 .extended_lut = "off";
defparam \Equal1~0 .lut_mask = 64'hFFFDFFFDFFFDFFFD;
defparam \Equal1~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal2~0 (
	.dataa(!A_mem_baddr_12),
	.datab(!A_mem_baddr_11),
	.datac(!A_mem_baddr_10),
	.datad(!A_mem_baddr_9),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal2),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal2~0 .extended_lut = "off";
defparam \Equal2~0 .lut_mask = 64'hFFFDFFFDFFFDFFFD;
defparam \Equal2~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal15~1 (
	.dataa(!A_mem_baddr_4),
	.datab(!A_mem_baddr_5),
	.datac(!A_mem_baddr_8),
	.datad(!Equal1),
	.datae(!Equal2),
	.dataf(!\Equal15~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal15),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal15~1 .extended_lut = "off";
defparam \Equal15~1 .lut_mask = 64'hFBFFFFFFFFFFFFFF;
defparam \Equal15~1 .shared_arith = "off";

cyclonev_lcell_comb \Equal14~0 (
	.dataa(!A_mem_baddr_4),
	.datab(!A_mem_baddr_7),
	.datac(!A_mem_baddr_6),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal14),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal14~0 .extended_lut = "off";
defparam \Equal14~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \Equal14~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal6~0 (
	.dataa(!A_mem_baddr_4),
	.datab(!A_mem_baddr_6),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal6),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal6~0 .extended_lut = "off";
defparam \Equal6~0 .lut_mask = 64'h7777777777777777;
defparam \Equal6~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal6~1 (
	.dataa(!A_mem_baddr_7),
	.datab(!A_mem_baddr_5),
	.datac(!A_mem_baddr_8),
	.datad(!Equal1),
	.datae(!Equal2),
	.dataf(!Equal6),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal61),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal6~1 .extended_lut = "off";
defparam \Equal6~1 .lut_mask = 64'hFEFFFFFFFFFFFFFF;
defparam \Equal6~1 .shared_arith = "off";

cyclonev_lcell_comb \always1~0 (
	.dataa(!A_mem_baddr_4),
	.datab(!A_mem_baddr_6),
	.datac(!A_mem_baddr_5),
	.datad(!A_mem_baddr_8),
	.datae(!Equal1),
	.dataf(!Equal2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(always1),
	.sumout(),
	.cout(),
	.shareout());
defparam \always1~0 .extended_lut = "off";
defparam \always1~0 .lut_mask = 64'hFFFBFFFFFFFFFFFF;
defparam \always1~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal16~0 (
	.dataa(!A_mem_baddr_4),
	.datab(!A_mem_baddr_5),
	.datac(!A_mem_baddr_8),
	.datad(!Equal1),
	.datae(!Equal2),
	.dataf(!\Equal15~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal16),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal16~0 .extended_lut = "off";
defparam \Equal16~0 .lut_mask = 64'hF7FFFFFFFFFFFFFF;
defparam \Equal16~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal2~1 (
	.dataa(!A_mem_baddr_5),
	.datab(!A_mem_baddr_8),
	.datac(!Equal1),
	.datad(!Equal2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal21),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal2~1 .extended_lut = "off";
defparam \Equal2~1 .lut_mask = 64'hEFFFEFFFEFFFEFFF;
defparam \Equal2~1 .shared_arith = "off";

cyclonev_lcell_comb \Equal2~2 (
	.dataa(!A_mem_baddr_7),
	.datab(!A_mem_baddr_6),
	.datac(!A_mem_baddr_5),
	.datad(!A_mem_baddr_8),
	.datae(!Equal1),
	.dataf(!Equal2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal22),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal2~2 .extended_lut = "off";
defparam \Equal2~2 .lut_mask = 64'hFFFEFFFFFFFFFFFF;
defparam \Equal2~2 .shared_arith = "off";

cyclonev_lcell_comb \always1~1 (
	.dataa(!A_mem_baddr_7),
	.datab(!A_mem_baddr_5),
	.datac(!A_mem_baddr_8),
	.datad(!Equal1),
	.datae(!Equal2),
	.dataf(!uav_read),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(always11),
	.sumout(),
	.cout(),
	.shareout());
defparam \always1~1 .extended_lut = "off";
defparam \always1~1 .lut_mask = 64'hFBFFFFFFFFFFFFFF;
defparam \always1~1 .shared_arith = "off";

cyclonev_lcell_comb \always1~2 (
	.dataa(!A_mem_baddr_7),
	.datab(!A_mem_baddr_6),
	.datac(!A_mem_baddr_5),
	.datad(!A_mem_baddr_8),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(always12),
	.sumout(),
	.cout(),
	.shareout());
defparam \always1~2 .extended_lut = "off";
defparam \always1~2 .lut_mask = 64'hFEFFFEFFFEFFFEFF;
defparam \always1~2 .shared_arith = "off";

cyclonev_lcell_comb \src_channel[2]~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\Equal15~2_combout ),
	.datad(!always11),
	.datae(!\src_channel[2]~0_combout ),
	.dataf(!\src_channel[2]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_channel_2),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_channel[2]~2 .extended_lut = "off";
defparam \src_channel[2]~2 .lut_mask = 64'hFFFFFFFFFFFFFFF0;
defparam \src_channel[2]~2 .shared_arith = "off";

cyclonev_lcell_comb \src_channel[2]~3 (
	.dataa(!A_mem_baddr_4),
	.datab(!A_mem_baddr_7),
	.datac(!A_mem_baddr_6),
	.datad(!A_mem_baddr_5),
	.datae(!\Equal2~3_combout ),
	.dataf(!uav_read),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_channel_21),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_channel[2]~3 .extended_lut = "off";
defparam \src_channel[2]~3 .lut_mask = 64'hFFB8FFFFFFFFFFFF;
defparam \src_channel[2]~3 .shared_arith = "off";

cyclonev_lcell_comb \Equal1~1 (
	.dataa(!A_mem_baddr_12),
	.datab(!A_mem_baddr_11),
	.datac(!A_mem_baddr_16),
	.datad(!A_mem_baddr_15),
	.datae(!A_mem_baddr_14),
	.dataf(!A_mem_baddr_13),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal11),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal1~1 .extended_lut = "off";
defparam \Equal1~1 .lut_mask = 64'hFFFFFFFFFFFFFFBF;
defparam \Equal1~1 .shared_arith = "off";

cyclonev_lcell_comb \always1~3 (
	.dataa(!A_mem_baddr_7),
	.datab(!always1),
	.datac(!uav_read),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(always13),
	.sumout(),
	.cout(),
	.shareout());
defparam \always1~3 .extended_lut = "off";
defparam \always1~3 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \always1~3 .shared_arith = "off";

cyclonev_lcell_comb \always1~4 (
	.dataa(!A_mem_baddr_4),
	.datab(!A_mem_baddr_6),
	.datac(!always11),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(always14),
	.sumout(),
	.cout(),
	.shareout());
defparam \always1~4 .extended_lut = "off";
defparam \always1~4 .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \always1~4 .shared_arith = "off";

cyclonev_lcell_comb \always1~5 (
	.dataa(!A_mem_baddr_4),
	.datab(!A_mem_baddr_6),
	.datac(!always11),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(always15),
	.sumout(),
	.cout(),
	.shareout());
defparam \always1~5 .extended_lut = "off";
defparam \always1~5 .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \always1~5 .shared_arith = "off";

cyclonev_lcell_comb \always1~6 (
	.dataa(!A_mem_baddr_4),
	.datab(!A_mem_baddr_6),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(always16),
	.sumout(),
	.cout(),
	.shareout());
defparam \always1~6 .extended_lut = "off";
defparam \always1~6 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \always1~6 .shared_arith = "off";

cyclonev_lcell_comb \always1~7 (
	.dataa(!A_mem_baddr_3),
	.datab(!A_mem_baddr_4),
	.datac(!Equal1),
	.datad(!Equal2),
	.datae(!uav_read),
	.dataf(!always12),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(always17),
	.sumout(),
	.cout(),
	.shareout());
defparam \always1~7 .extended_lut = "off";
defparam \always1~7 .lut_mask = 64'hEFFFFFFFFFFFFFFF;
defparam \always1~7 .shared_arith = "off";

cyclonev_lcell_comb \always1~9 (
	.dataa(!A_mem_baddr_5),
	.datab(!A_mem_baddr_8),
	.datac(!Equal1),
	.datad(!Equal2),
	.datae(!uav_read),
	.dataf(!\always1~8_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(always18),
	.sumout(),
	.cout(),
	.shareout());
defparam \always1~9 .extended_lut = "off";
defparam \always1~9 .lut_mask = 64'hDFFFFFFFFFFFFFFF;
defparam \always1~9 .shared_arith = "off";

cyclonev_lcell_comb \always1~11 (
	.dataa(!A_mem_baddr_5),
	.datab(!A_mem_baddr_8),
	.datac(!Equal1),
	.datad(!Equal2),
	.datae(!uav_read),
	.dataf(!\always1~10_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(always19),
	.sumout(),
	.cout(),
	.shareout());
defparam \always1~11 .extended_lut = "off";
defparam \always1~11 .lut_mask = 64'hDFFFFFFFFFFFFFFF;
defparam \always1~11 .shared_arith = "off";

cyclonev_lcell_comb \always1~12 (
	.dataa(!A_mem_baddr_5),
	.datab(!A_mem_baddr_8),
	.datac(!Equal1),
	.datad(!Equal2),
	.datae(!uav_read),
	.dataf(!\always1~8_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(always110),
	.sumout(),
	.cout(),
	.shareout());
defparam \always1~12 .extended_lut = "off";
defparam \always1~12 .lut_mask = 64'hEFFFFFFFFFFFFFFF;
defparam \always1~12 .shared_arith = "off";

cyclonev_lcell_comb \always1~13 (
	.dataa(!Equal1),
	.datab(!Equal2),
	.datac(!always12),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(always111),
	.sumout(),
	.cout(),
	.shareout());
defparam \always1~13 .extended_lut = "off";
defparam \always1~13 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \always1~13 .shared_arith = "off";

cyclonev_lcell_comb \Equal15~0 (
	.dataa(!A_mem_baddr_7),
	.datab(!A_mem_baddr_6),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal15~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal15~0 .extended_lut = "off";
defparam \Equal15~0 .lut_mask = 64'h7777777777777777;
defparam \Equal15~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal15~2 (
	.dataa(!A_mem_baddr_5),
	.datab(!A_mem_baddr_8),
	.datac(!Equal1),
	.datad(!Equal2),
	.datae(!\Equal15~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal15~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal15~2 .extended_lut = "off";
defparam \Equal15~2 .lut_mask = 64'hDFFFFFFFDFFFFFFF;
defparam \Equal15~2 .shared_arith = "off";

cyclonev_lcell_comb \src_channel[2]~0 (
	.dataa(gnd),
	.datab(!A_mem_baddr_5),
	.datac(!A_mem_baddr_8),
	.datad(!Equal1),
	.datae(!Equal2),
	.dataf(!Equal6),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_channel[2]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_channel[2]~0 .extended_lut = "off";
defparam \src_channel[2]~0 .lut_mask = 64'hFCFFFFFFFFFFFFFF;
defparam \src_channel[2]~0 .shared_arith = "off";

cyclonev_lcell_comb \src_channel[2]~1 (
	.dataa(!A_mem_baddr_3),
	.datab(!A_mem_baddr_4),
	.datac(!Equal1),
	.datad(!Equal2),
	.datae(!uav_read),
	.dataf(!always12),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_channel[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_channel[2]~1 .extended_lut = "off";
defparam \src_channel[2]~1 .lut_mask = 64'hDFFFFFFFFFFFFFFF;
defparam \src_channel[2]~1 .shared_arith = "off";

cyclonev_lcell_comb \Equal2~3 (
	.dataa(!A_mem_baddr_8),
	.datab(!Equal1),
	.datac(!Equal2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal2~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal2~3 .extended_lut = "off";
defparam \Equal2~3 .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \Equal2~3 .shared_arith = "off";

cyclonev_lcell_comb \always1~8 (
	.dataa(!A_mem_baddr_4),
	.datab(!A_mem_baddr_7),
	.datac(!A_mem_baddr_6),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always1~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always1~8 .extended_lut = "off";
defparam \always1~8 .lut_mask = 64'hF7F7F7F7F7F7F7F7;
defparam \always1~8 .shared_arith = "off";

cyclonev_lcell_comb \always1~10 (
	.dataa(!A_mem_baddr_4),
	.datab(!A_mem_baddr_7),
	.datac(!A_mem_baddr_6),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always1~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always1~10 .extended_lut = "off";
defparam \always1~10 .lut_mask = 64'hFBFBFBFBFBFBFBFB;
defparam \always1~10 .shared_arith = "off";

endmodule

module first_nios2_system_first_nios2_system_mm_interconnect_0_router_001 (
	ic_fill_tag_5,
	ic_fill_tag_4,
	ic_fill_tag_3,
	ic_fill_tag_2,
	ic_fill_tag_1,
	ic_fill_tag_0,
	Equal1)/* synthesis synthesis_greybox=1 */;
input 	ic_fill_tag_5;
input 	ic_fill_tag_4;
input 	ic_fill_tag_3;
input 	ic_fill_tag_2;
input 	ic_fill_tag_1;
input 	ic_fill_tag_0;
output 	Equal1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \Equal1~0 (
	.dataa(!ic_fill_tag_5),
	.datab(!ic_fill_tag_4),
	.datac(!ic_fill_tag_3),
	.datad(!ic_fill_tag_2),
	.datae(!ic_fill_tag_1),
	.dataf(!ic_fill_tag_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal1),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal1~0 .extended_lut = "off";
defparam \Equal1~0 .lut_mask = 64'hFFFFFFFDFFFFFFFF;
defparam \Equal1~0 .shared_arith = "off";

endmodule

module first_nios2_system_first_nios2_system_mm_interconnect_0_rsp_demux_002 (
	read_latency_shift_reg_0,
	mem_74_0,
	mem_56_0,
	src0_valid,
	src1_valid)/* synthesis synthesis_greybox=1 */;
input 	read_latency_shift_reg_0;
input 	mem_74_0;
input 	mem_56_0;
output 	src0_valid;
output 	src1_valid;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \src0_valid~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_74_0),
	.datac(!mem_56_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src0_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src0_valid~0 .extended_lut = "off";
defparam \src0_valid~0 .lut_mask = 64'hFDFDFDFDFDFDFDFD;
defparam \src0_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \src1_valid~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_74_0),
	.datac(!mem_56_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src1_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src1_valid~0 .extended_lut = "off";
defparam \src1_valid~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \src1_valid~0 .shared_arith = "off";

endmodule

module first_nios2_system_first_nios2_system_mm_interconnect_0_rsp_demux_002_1 (
	read_latency_shift_reg_0,
	mem_74_0,
	mem_56_0,
	src0_valid,
	src1_valid)/* synthesis synthesis_greybox=1 */;
input 	read_latency_shift_reg_0;
input 	mem_74_0;
input 	mem_56_0;
output 	src0_valid;
output 	src1_valid;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \src0_valid~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_74_0),
	.datac(!mem_56_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src0_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src0_valid~0 .extended_lut = "off";
defparam \src0_valid~0 .lut_mask = 64'hFDFDFDFDFDFDFDFD;
defparam \src0_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \src1_valid~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_74_0),
	.datac(!mem_56_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src1_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src1_valid~0 .extended_lut = "off";
defparam \src1_valid~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \src1_valid~0 .shared_arith = "off";

endmodule

module first_nios2_system_first_nios2_system_mm_interconnect_0_rsp_mux (
	av_readdata_pre_0,
	q_a_0,
	av_readdata_pre_01,
	av_readdata_pre_02,
	av_readdata_pre_03,
	av_readdata_pre_04,
	av_readdata_pre_05,
	av_readdata_pre_06,
	av_readdata_pre_1,
	q_a_1,
	av_readdata_pre_11,
	av_readdata_pre_12,
	av_readdata_pre_13,
	av_readdata_pre_2,
	q_a_2,
	av_readdata_pre_21,
	av_readdata_pre_22,
	av_readdata_pre_23,
	q_a_3,
	av_readdata_pre_3,
	av_readdata_pre_31,
	av_readdata_pre_32,
	av_readdata_pre_33,
	av_readdata_pre_4,
	av_readdata_pre_41,
	q_a_4,
	av_readdata_pre_42,
	av_readdata_pre_43,
	av_readdata_pre_5,
	q_a_5,
	av_readdata_pre_51,
	av_readdata_pre_52,
	av_readdata_pre_53,
	q_a_6,
	av_readdata_pre_6,
	av_readdata_pre_61,
	av_readdata_pre_62,
	av_readdata_pre_63,
	q_a_7,
	av_readdata_pre_7,
	av_readdata_pre_71,
	av_readdata_pre_221,
	q_a_22,
	q_a_23,
	q_a_24,
	q_a_25,
	q_a_31,
	q_a_21,
	av_readdata_pre_211,
	q_a_11,
	q_a_28,
	q_a_10,
	q_a_27,
	q_a_8,
	q_a_9,
	q_a_26,
	av_readdata_pre_20,
	q_a_20,
	av_readdata_pre_19,
	q_a_19,
	q_a_17,
	av_readdata_pre_17,
	q_a_30,
	q_a_18,
	av_readdata_pre_18,
	q_a_16,
	av_readdata_pre_16,
	q_a_15,
	q_a_12,
	q_a_13,
	q_a_14,
	q_a_29,
	read_latency_shift_reg_0,
	read_latency_shift_reg_01,
	read_latency_shift_reg_02,
	read_latency_shift_reg_03,
	read_latency_shift_reg_04,
	read_latency_shift_reg_05,
	read_latency_shift_reg_06,
	WideOr11,
	read_latency_shift_reg_07,
	read_latency_shift_reg_08,
	read_latency_shift_reg_09,
	read_latency_shift_reg_010,
	read_latency_shift_reg_011,
	WideOr12,
	read_latency_shift_reg_012,
	src0_valid,
	src0_valid1,
	read_latency_shift_reg_013,
	read_latency_shift_reg_014,
	read_latency_shift_reg_015,
	read_latency_shift_reg_016,
	WideOr13,
	WideOr14,
	av_readdata_pre_07,
	av_readdata_pre_08,
	av_readdata_pre_09,
	av_readdata_pre_010,
	av_readdata_pre_011,
	av_readdata_pre_012,
	av_readdata_pre_013,
	av_readdata_pre_014,
	av_readdata_pre_015,
	av_readdata_pre_016,
	src_data_0,
	av_readdata_pre_14,
	av_readdata_pre_15,
	av_readdata_pre_110,
	av_readdata_pre_111,
	av_readdata_pre_30,
	src_payload,
	av_readdata_pre_112,
	av_readdata_pre_113,
	av_readdata_pre_114,
	av_readdata_pre_115,
	src_data_1,
	av_readdata_pre_24,
	av_readdata_pre_25,
	av_readdata_pre_26,
	av_readdata_pre_27,
	av_readdata_pre_28,
	av_readdata_pre_29,
	av_readdata_pre_210,
	av_readdata_pre_212,
	src_data_2,
	av_readdata_pre_34,
	av_readdata_pre_35,
	av_readdata_pre_36,
	av_readdata_pre_37,
	av_readdata_pre_38,
	av_readdata_pre_39,
	av_readdata_pre_310,
	av_readdata_pre_311,
	src_data_3,
	av_readdata_pre_44,
	av_readdata_pre_45,
	av_readdata_pre_46,
	av_readdata_pre_47,
	av_readdata_pre_48,
	av_readdata_pre_49,
	src_payload1,
	av_readdata_pre_54,
	av_readdata_pre_55,
	av_readdata_pre_56,
	av_readdata_pre_57,
	av_readdata_pre_58,
	av_readdata_pre_59,
	src_payload2,
	av_readdata_pre_64,
	av_readdata_pre_65,
	av_readdata_pre_66,
	av_readdata_pre_67,
	src_payload3,
	av_readdata_pre_72,
	av_readdata_pre_73,
	src_payload4,
	av_readdata_pre_222,
	src_payload5,
	av_readdata_pre_231,
	src_payload6,
	av_readdata_pre_241,
	src_payload7,
	av_readdata_pre_251,
	src_payload8,
	av_readdata_pre_312,
	src_payload9,
	av_readdata_pre_213,
	src_payload10,
	src_payload11,
	av_readdata_pre_116,
	av_readdata_pre_117,
	src_payload12,
	src_payload13,
	av_readdata_pre_281,
	src_payload14,
	av_readdata_pre_10,
	av_readdata_pre_101,
	av_readdata_pre_102,
	src_payload15,
	src_payload16,
	av_readdata_pre_271,
	src_payload17,
	av_readdata_pre_8,
	av_readdata_pre_81,
	av_readdata_pre_82,
	src_payload18,
	src_payload19,
	av_readdata_pre_9,
	av_readdata_pre_91,
	av_readdata_pre_92,
	src_payload20,
	src_payload21,
	av_readdata_pre_261,
	src_payload22,
	av_readdata_pre_201,
	src_payload23,
	av_readdata_pre_191,
	src_payload24,
	av_readdata_pre_171,
	src_payload25,
	src_payload26,
	av_readdata_pre_301,
	src_payload27,
	av_readdata_pre_181,
	src_payload28,
	src_payload29,
	av_readdata_pre_161,
	src_payload30,
	src_payload31,
	av_readdata_pre_151,
	av_readdata_pre_152,
	av_readdata_pre_153,
	src_payload32,
	src_payload33,
	av_readdata_pre_121,
	av_readdata_pre_122,
	av_readdata_pre_123,
	src_payload34,
	src_payload35,
	av_readdata_pre_131,
	av_readdata_pre_132,
	av_readdata_pre_133,
	src_payload36,
	src_payload37,
	av_readdata_pre_141,
	av_readdata_pre_142,
	av_readdata_pre_143,
	src_payload38,
	src_payload39,
	av_readdata_pre_291,
	src_payload40)/* synthesis synthesis_greybox=1 */;
input 	av_readdata_pre_0;
input 	q_a_0;
input 	av_readdata_pre_01;
input 	av_readdata_pre_02;
input 	av_readdata_pre_03;
input 	av_readdata_pre_04;
input 	av_readdata_pre_05;
input 	av_readdata_pre_06;
input 	av_readdata_pre_1;
input 	q_a_1;
input 	av_readdata_pre_11;
input 	av_readdata_pre_12;
input 	av_readdata_pre_13;
input 	av_readdata_pre_2;
input 	q_a_2;
input 	av_readdata_pre_21;
input 	av_readdata_pre_22;
input 	av_readdata_pre_23;
input 	q_a_3;
input 	av_readdata_pre_3;
input 	av_readdata_pre_31;
input 	av_readdata_pre_32;
input 	av_readdata_pre_33;
input 	av_readdata_pre_4;
input 	av_readdata_pre_41;
input 	q_a_4;
input 	av_readdata_pre_42;
input 	av_readdata_pre_43;
input 	av_readdata_pre_5;
input 	q_a_5;
input 	av_readdata_pre_51;
input 	av_readdata_pre_52;
input 	av_readdata_pre_53;
input 	q_a_6;
input 	av_readdata_pre_6;
input 	av_readdata_pre_61;
input 	av_readdata_pre_62;
input 	av_readdata_pre_63;
input 	q_a_7;
input 	av_readdata_pre_7;
input 	av_readdata_pre_71;
input 	av_readdata_pre_221;
input 	q_a_22;
input 	q_a_23;
input 	q_a_24;
input 	q_a_25;
input 	q_a_31;
input 	q_a_21;
input 	av_readdata_pre_211;
input 	q_a_11;
input 	q_a_28;
input 	q_a_10;
input 	q_a_27;
input 	q_a_8;
input 	q_a_9;
input 	q_a_26;
input 	av_readdata_pre_20;
input 	q_a_20;
input 	av_readdata_pre_19;
input 	q_a_19;
input 	q_a_17;
input 	av_readdata_pre_17;
input 	q_a_30;
input 	q_a_18;
input 	av_readdata_pre_18;
input 	q_a_16;
input 	av_readdata_pre_16;
input 	q_a_15;
input 	q_a_12;
input 	q_a_13;
input 	q_a_14;
input 	q_a_29;
input 	read_latency_shift_reg_0;
input 	read_latency_shift_reg_01;
input 	read_latency_shift_reg_02;
input 	read_latency_shift_reg_03;
input 	read_latency_shift_reg_04;
input 	read_latency_shift_reg_05;
input 	read_latency_shift_reg_06;
output 	WideOr11;
input 	read_latency_shift_reg_07;
input 	read_latency_shift_reg_08;
input 	read_latency_shift_reg_09;
input 	read_latency_shift_reg_010;
input 	read_latency_shift_reg_011;
output 	WideOr12;
input 	read_latency_shift_reg_012;
input 	src0_valid;
input 	src0_valid1;
input 	read_latency_shift_reg_013;
input 	read_latency_shift_reg_014;
input 	read_latency_shift_reg_015;
input 	read_latency_shift_reg_016;
output 	WideOr13;
output 	WideOr14;
input 	av_readdata_pre_07;
input 	av_readdata_pre_08;
input 	av_readdata_pre_09;
input 	av_readdata_pre_010;
input 	av_readdata_pre_011;
input 	av_readdata_pre_012;
input 	av_readdata_pre_013;
input 	av_readdata_pre_014;
input 	av_readdata_pre_015;
input 	av_readdata_pre_016;
output 	src_data_0;
input 	av_readdata_pre_14;
input 	av_readdata_pre_15;
input 	av_readdata_pre_110;
input 	av_readdata_pre_111;
input 	av_readdata_pre_30;
output 	src_payload;
input 	av_readdata_pre_112;
input 	av_readdata_pre_113;
input 	av_readdata_pre_114;
input 	av_readdata_pre_115;
output 	src_data_1;
input 	av_readdata_pre_24;
input 	av_readdata_pre_25;
input 	av_readdata_pre_26;
input 	av_readdata_pre_27;
input 	av_readdata_pre_28;
input 	av_readdata_pre_29;
input 	av_readdata_pre_210;
input 	av_readdata_pre_212;
output 	src_data_2;
input 	av_readdata_pre_34;
input 	av_readdata_pre_35;
input 	av_readdata_pre_36;
input 	av_readdata_pre_37;
input 	av_readdata_pre_38;
input 	av_readdata_pre_39;
input 	av_readdata_pre_310;
input 	av_readdata_pre_311;
output 	src_data_3;
input 	av_readdata_pre_44;
input 	av_readdata_pre_45;
input 	av_readdata_pre_46;
input 	av_readdata_pre_47;
input 	av_readdata_pre_48;
input 	av_readdata_pre_49;
output 	src_payload1;
input 	av_readdata_pre_54;
input 	av_readdata_pre_55;
input 	av_readdata_pre_56;
input 	av_readdata_pre_57;
input 	av_readdata_pre_58;
input 	av_readdata_pre_59;
output 	src_payload2;
input 	av_readdata_pre_64;
input 	av_readdata_pre_65;
input 	av_readdata_pre_66;
input 	av_readdata_pre_67;
output 	src_payload3;
input 	av_readdata_pre_72;
input 	av_readdata_pre_73;
output 	src_payload4;
input 	av_readdata_pre_222;
output 	src_payload5;
input 	av_readdata_pre_231;
output 	src_payload6;
input 	av_readdata_pre_241;
output 	src_payload7;
input 	av_readdata_pre_251;
output 	src_payload8;
input 	av_readdata_pre_312;
output 	src_payload9;
input 	av_readdata_pre_213;
output 	src_payload10;
output 	src_payload11;
input 	av_readdata_pre_116;
input 	av_readdata_pre_117;
output 	src_payload12;
output 	src_payload13;
input 	av_readdata_pre_281;
output 	src_payload14;
input 	av_readdata_pre_10;
input 	av_readdata_pre_101;
input 	av_readdata_pre_102;
output 	src_payload15;
output 	src_payload16;
input 	av_readdata_pre_271;
output 	src_payload17;
input 	av_readdata_pre_8;
input 	av_readdata_pre_81;
input 	av_readdata_pre_82;
output 	src_payload18;
output 	src_payload19;
input 	av_readdata_pre_9;
input 	av_readdata_pre_91;
input 	av_readdata_pre_92;
output 	src_payload20;
output 	src_payload21;
input 	av_readdata_pre_261;
output 	src_payload22;
input 	av_readdata_pre_201;
output 	src_payload23;
input 	av_readdata_pre_191;
output 	src_payload24;
input 	av_readdata_pre_171;
output 	src_payload25;
output 	src_payload26;
input 	av_readdata_pre_301;
output 	src_payload27;
input 	av_readdata_pre_181;
output 	src_payload28;
output 	src_payload29;
input 	av_readdata_pre_161;
output 	src_payload30;
output 	src_payload31;
input 	av_readdata_pre_151;
input 	av_readdata_pre_152;
input 	av_readdata_pre_153;
output 	src_payload32;
output 	src_payload33;
input 	av_readdata_pre_121;
input 	av_readdata_pre_122;
input 	av_readdata_pre_123;
output 	src_payload34;
output 	src_payload35;
input 	av_readdata_pre_131;
input 	av_readdata_pre_132;
input 	av_readdata_pre_133;
output 	src_payload36;
output 	src_payload37;
input 	av_readdata_pre_141;
input 	av_readdata_pre_142;
input 	av_readdata_pre_143;
output 	src_payload38;
output 	src_payload39;
input 	av_readdata_pre_291;
output 	src_payload40;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \WideOr1~2_combout ;
wire \src_data[0]~0_combout ;
wire \src_data[0]~3_combout ;
wire \src_data[0]~4_combout ;
wire \src_data[0]~5_combout ;
wire \src_data[0]~18_combout ;
wire \src_data[0]~1_combout ;
wire \src_data[0]~2_combout ;
wire \src_data[0]~19_combout ;
wire \src_data[1]~6_combout ;
wire \src_data[1]~7_combout ;
wire \src_data[1]~20_combout ;
wire \src_data[1]~8_combout ;
wire \src_data[1]~21_combout ;
wire \src_data[2]~9_combout ;
wire \src_data[2]~10_combout ;
wire \src_data[2]~22_combout ;
wire \src_data[2]~11_combout ;
wire \src_data[2]~23_combout ;
wire \src_data[3]~12_combout ;
wire \src_data[3]~13_combout ;
wire \src_data[3]~14_combout ;
wire \src_data[3]~15_combout ;
wire \src_data[3]~16_combout ;
wire \src_data[3]~17_combout ;
wire \src_payload~1_combout ;
wire \src_payload~2_combout ;
wire \src_payload~52_combout ;
wire \src_payload~53_combout ;
wire \src_payload~4_combout ;
wire \src_payload~5_combout ;
wire \src_payload~6_combout ;
wire \src_payload~54_combout ;
wire \src_payload~8_combout ;
wire \src_payload~9_combout ;
wire \src_payload~10_combout ;
wire \src_payload~11_combout ;
wire \src_payload~13_combout ;
wire \src_payload~14_combout ;


cyclonev_lcell_comb \WideOr1~0 (
	.dataa(!read_latency_shift_reg_02),
	.datab(!read_latency_shift_reg_03),
	.datac(!read_latency_shift_reg_04),
	.datad(!read_latency_shift_reg_05),
	.datae(!read_latency_shift_reg_06),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr11),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr1~0 .extended_lut = "off";
defparam \WideOr1~0 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \WideOr1~0 .shared_arith = "off";

cyclonev_lcell_comb \WideOr1~1 (
	.dataa(!read_latency_shift_reg_07),
	.datab(!read_latency_shift_reg_08),
	.datac(!read_latency_shift_reg_09),
	.datad(!read_latency_shift_reg_010),
	.datae(!read_latency_shift_reg_011),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr12),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr1~1 .extended_lut = "off";
defparam \WideOr1~1 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \WideOr1~1 .shared_arith = "off";

cyclonev_lcell_comb \WideOr1~3 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!read_latency_shift_reg_012),
	.datac(!src0_valid),
	.datad(!src0_valid1),
	.datae(!\WideOr1~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr13),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr1~3 .extended_lut = "off";
defparam \WideOr1~3 .lut_mask = 64'hFFFEFFFFFFFEFFFF;
defparam \WideOr1~3 .shared_arith = "off";

cyclonev_lcell_comb WideOr1(
	.dataa(!read_latency_shift_reg_01),
	.datab(!WideOr11),
	.datac(!WideOr12),
	.datad(!WideOr13),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr14),
	.sumout(),
	.cout(),
	.shareout());
defparam WideOr1.extended_lut = "off";
defparam WideOr1.lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam WideOr1.shared_arith = "off";

cyclonev_lcell_comb \src_data[0] (
	.dataa(!\src_data[0]~0_combout ),
	.datab(!src0_valid1),
	.datac(!q_a_0),
	.datad(!\src_data[0]~5_combout ),
	.datae(!\src_data[0]~18_combout ),
	.dataf(!\src_data[0]~19_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[0] .extended_lut = "off";
defparam \src_data[0] .lut_mask = 64'hFFFFFFFFFFFFFFBF;
defparam \src_data[0] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~0 (
	.dataa(!read_latency_shift_reg_014),
	.datab(!av_readdata_pre_30),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~0 .extended_lut = "off";
defparam \src_payload~0 .lut_mask = 64'h7777777777777777;
defparam \src_payload~0 .shared_arith = "off";

cyclonev_lcell_comb \src_data[1] (
	.dataa(!src0_valid1),
	.datab(!q_a_1),
	.datac(!\src_data[1]~6_combout ),
	.datad(!\src_data[1]~7_combout ),
	.datae(!\src_data[1]~20_combout ),
	.dataf(!\src_data[1]~21_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[1] .extended_lut = "off";
defparam \src_data[1] .lut_mask = 64'hFFFFFFFFFFFFF7FF;
defparam \src_data[1] .shared_arith = "off";

cyclonev_lcell_comb \src_data[2] (
	.dataa(!src0_valid1),
	.datab(!q_a_2),
	.datac(!\src_data[2]~9_combout ),
	.datad(!\src_data[2]~10_combout ),
	.datae(!\src_data[2]~22_combout ),
	.dataf(!\src_data[2]~23_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_2),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[2] .extended_lut = "off";
defparam \src_data[2] .lut_mask = 64'hFFFFFFFFFFFFF7FF;
defparam \src_data[2] .shared_arith = "off";

cyclonev_lcell_comb \src_data[3] (
	.dataa(!read_latency_shift_reg_08),
	.datab(!src0_valid1),
	.datac(!q_a_3),
	.datad(!av_readdata_pre_34),
	.datae(!\src_data[3]~17_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_3),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[3] .extended_lut = "off";
defparam \src_data[3] .lut_mask = 64'hFFFF7FFFFFFF7FFF;
defparam \src_data[3] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~3 (
	.dataa(!\src_payload~1_combout ),
	.datab(!\src_payload~2_combout ),
	.datac(!src0_valid1),
	.datad(!q_a_4),
	.datae(!\src_payload~52_combout ),
	.dataf(!\src_payload~53_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~3 .extended_lut = "off";
defparam \src_payload~3 .lut_mask = 64'hFFFFFFFFFFFFBFFF;
defparam \src_payload~3 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~7 (
	.dataa(!\src_payload~6_combout ),
	.datab(!src0_valid1),
	.datac(!q_a_5),
	.datad(!read_latency_shift_reg_07),
	.datae(!av_readdata_pre_55),
	.dataf(!\src_payload~54_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload2),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~7 .extended_lut = "off";
defparam \src_payload~7 .lut_mask = 64'hFFFFFFFFBFFFFFFF;
defparam \src_payload~7 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~12 (
	.dataa(!read_latency_shift_reg_07),
	.datab(!src0_valid1),
	.datac(!q_a_6),
	.datad(!av_readdata_pre_64),
	.datae(!\src_payload~11_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload3),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~12 .extended_lut = "off";
defparam \src_payload~12 .lut_mask = 64'hFFFF7FFFFFFF7FFF;
defparam \src_payload~12 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~15 (
	.dataa(!src0_valid1),
	.datab(!q_a_7),
	.datac(!\src_payload~13_combout ),
	.datad(!\src_payload~14_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload4),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~15 .extended_lut = "off";
defparam \src_payload~15 .lut_mask = 64'hF7FFF7FFF7FFF7FF;
defparam \src_payload~15 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~16 (
	.dataa(!read_latency_shift_reg_013),
	.datab(!src0_valid),
	.datac(!src0_valid1),
	.datad(!av_readdata_pre_221),
	.datae(!av_readdata_pre_222),
	.dataf(!q_a_22),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload5),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~16 .extended_lut = "off";
defparam \src_payload~16 .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \src_payload~16 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~17 (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!av_readdata_pre_231),
	.datad(!q_a_23),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload6),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~17 .extended_lut = "off";
defparam \src_payload~17 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_payload~17 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~18 (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!av_readdata_pre_241),
	.datad(!q_a_24),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload7),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~18 .extended_lut = "off";
defparam \src_payload~18 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_payload~18 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~19 (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!src_payload),
	.datad(!av_readdata_pre_251),
	.datae(!q_a_25),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload8),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~19 .extended_lut = "off";
defparam \src_payload~19 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \src_payload~19 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~20 (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!av_readdata_pre_312),
	.datad(!q_a_31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload9),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~20 .extended_lut = "off";
defparam \src_payload~20 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_payload~20 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~21 (
	.dataa(!read_latency_shift_reg_013),
	.datab(!src_payload),
	.datac(!av_readdata_pre_211),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload10),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~21 .extended_lut = "off";
defparam \src_payload~21 .lut_mask = 64'hFEFEFEFEFEFEFEFE;
defparam \src_payload~21 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~22 (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!av_readdata_pre_213),
	.datad(!q_a_21),
	.datae(!src_payload10),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload11),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~22 .extended_lut = "off";
defparam \src_payload~22 .lut_mask = 64'hFFFF7FFFFFFF7FFF;
defparam \src_payload~22 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~23 (
	.dataa(!read_latency_shift_reg_015),
	.datab(!src_payload),
	.datac(!av_readdata_pre_117),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload12),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~23 .extended_lut = "off";
defparam \src_payload~23 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \src_payload~23 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~24 (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!av_readdata_pre_116),
	.datad(!q_a_11),
	.datae(!src_payload12),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload13),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~24 .extended_lut = "off";
defparam \src_payload~24 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \src_payload~24 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~25 (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!src_payload),
	.datad(!av_readdata_pre_281),
	.datae(!q_a_28),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload14),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~25 .extended_lut = "off";
defparam \src_payload~25 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \src_payload~25 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~26 (
	.dataa(!read_latency_shift_reg_013),
	.datab(!read_latency_shift_reg_015),
	.datac(!av_readdata_pre_101),
	.datad(!av_readdata_pre_102),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload15),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~26 .extended_lut = "off";
defparam \src_payload~26 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_payload~26 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~27 (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!av_readdata_pre_10),
	.datad(!q_a_10),
	.datae(!src_payload15),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload16),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~27 .extended_lut = "off";
defparam \src_payload~27 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \src_payload~27 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~28 (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!src_payload),
	.datad(!av_readdata_pre_271),
	.datae(!q_a_27),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload17),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~28 .extended_lut = "off";
defparam \src_payload~28 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \src_payload~28 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~29 (
	.dataa(!read_latency_shift_reg_013),
	.datab(!read_latency_shift_reg_015),
	.datac(!av_readdata_pre_81),
	.datad(!av_readdata_pre_82),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload18),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~29 .extended_lut = "off";
defparam \src_payload~29 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_payload~29 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~30 (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!av_readdata_pre_8),
	.datad(!q_a_8),
	.datae(!src_payload18),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload19),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~30 .extended_lut = "off";
defparam \src_payload~30 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \src_payload~30 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~31 (
	.dataa(!read_latency_shift_reg_013),
	.datab(!read_latency_shift_reg_015),
	.datac(!av_readdata_pre_91),
	.datad(!av_readdata_pre_92),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload20),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~31 .extended_lut = "off";
defparam \src_payload~31 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_payload~31 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~32 (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!av_readdata_pre_9),
	.datad(!q_a_9),
	.datae(!src_payload20),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload21),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~32 .extended_lut = "off";
defparam \src_payload~32 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \src_payload~32 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~33 (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!av_readdata_pre_261),
	.datad(!q_a_26),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload22),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~33 .extended_lut = "off";
defparam \src_payload~33 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_payload~33 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~34 (
	.dataa(!read_latency_shift_reg_013),
	.datab(!src0_valid),
	.datac(!src0_valid1),
	.datad(!av_readdata_pre_20),
	.datae(!av_readdata_pre_201),
	.dataf(!q_a_20),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload23),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~34 .extended_lut = "off";
defparam \src_payload~34 .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \src_payload~34 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~35 (
	.dataa(!read_latency_shift_reg_013),
	.datab(!src0_valid),
	.datac(!src0_valid1),
	.datad(!av_readdata_pre_19),
	.datae(!av_readdata_pre_191),
	.dataf(!q_a_19),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload24),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~35 .extended_lut = "off";
defparam \src_payload~35 .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \src_payload~35 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~36 (
	.dataa(!read_latency_shift_reg_013),
	.datab(!src_payload),
	.datac(!av_readdata_pre_17),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload25),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~36 .extended_lut = "off";
defparam \src_payload~36 .lut_mask = 64'hFEFEFEFEFEFEFEFE;
defparam \src_payload~36 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~37 (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!av_readdata_pre_171),
	.datad(!q_a_17),
	.datae(!src_payload25),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload26),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~37 .extended_lut = "off";
defparam \src_payload~37 .lut_mask = 64'hFFFF7FFFFFFF7FFF;
defparam \src_payload~37 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~38 (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!src_payload),
	.datad(!av_readdata_pre_301),
	.datae(!q_a_30),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload27),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~38 .extended_lut = "off";
defparam \src_payload~38 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \src_payload~38 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~39 (
	.dataa(!read_latency_shift_reg_013),
	.datab(!src_payload),
	.datac(!av_readdata_pre_18),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload28),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~39 .extended_lut = "off";
defparam \src_payload~39 .lut_mask = 64'hFEFEFEFEFEFEFEFE;
defparam \src_payload~39 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~40 (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!av_readdata_pre_181),
	.datad(!q_a_18),
	.datae(!src_payload28),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload29),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~40 .extended_lut = "off";
defparam \src_payload~40 .lut_mask = 64'hFFFF7FFFFFFF7FFF;
defparam \src_payload~40 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~41 (
	.dataa(!read_latency_shift_reg_013),
	.datab(!src_payload),
	.datac(!av_readdata_pre_16),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload30),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~41 .extended_lut = "off";
defparam \src_payload~41 .lut_mask = 64'hFEFEFEFEFEFEFEFE;
defparam \src_payload~41 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~42 (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!av_readdata_pre_161),
	.datad(!q_a_16),
	.datae(!src_payload30),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload31),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~42 .extended_lut = "off";
defparam \src_payload~42 .lut_mask = 64'hFFFF7FFFFFFF7FFF;
defparam \src_payload~42 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~43 (
	.dataa(!read_latency_shift_reg_013),
	.datab(!read_latency_shift_reg_015),
	.datac(!av_readdata_pre_152),
	.datad(!av_readdata_pre_153),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload32),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~43 .extended_lut = "off";
defparam \src_payload~43 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_payload~43 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~44 (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!av_readdata_pre_151),
	.datad(!q_a_15),
	.datae(!src_payload32),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload33),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~44 .extended_lut = "off";
defparam \src_payload~44 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \src_payload~44 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~45 (
	.dataa(!read_latency_shift_reg_013),
	.datab(!read_latency_shift_reg_015),
	.datac(!src_payload),
	.datad(!av_readdata_pre_122),
	.datae(!av_readdata_pre_123),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload34),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~45 .extended_lut = "off";
defparam \src_payload~45 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \src_payload~45 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~46 (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!av_readdata_pre_121),
	.datad(!q_a_12),
	.datae(!src_payload34),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload35),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~46 .extended_lut = "off";
defparam \src_payload~46 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \src_payload~46 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~47 (
	.dataa(!read_latency_shift_reg_013),
	.datab(!read_latency_shift_reg_015),
	.datac(!av_readdata_pre_132),
	.datad(!av_readdata_pre_133),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload36),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~47 .extended_lut = "off";
defparam \src_payload~47 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_payload~47 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~48 (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!av_readdata_pre_131),
	.datad(!q_a_13),
	.datae(!src_payload36),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload37),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~48 .extended_lut = "off";
defparam \src_payload~48 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \src_payload~48 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~49 (
	.dataa(!read_latency_shift_reg_013),
	.datab(!read_latency_shift_reg_015),
	.datac(!src_payload),
	.datad(!av_readdata_pre_142),
	.datae(!av_readdata_pre_143),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload38),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~49 .extended_lut = "off";
defparam \src_payload~49 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \src_payload~49 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~50 (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!av_readdata_pre_141),
	.datad(!q_a_14),
	.datae(!src_payload38),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload39),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~50 .extended_lut = "off";
defparam \src_payload~50 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \src_payload~50 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~51 (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!av_readdata_pre_291),
	.datad(!q_a_29),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload40),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~51 .extended_lut = "off";
defparam \src_payload~51 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_payload~51 .shared_arith = "off";

cyclonev_lcell_comb \WideOr1~2 (
	.dataa(!read_latency_shift_reg_013),
	.datab(!read_latency_shift_reg_014),
	.datac(!read_latency_shift_reg_015),
	.datad(!read_latency_shift_reg_016),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr1~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr1~2 .extended_lut = "off";
defparam \WideOr1~2 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \WideOr1~2 .shared_arith = "off";

cyclonev_lcell_comb \src_data[0]~0 (
	.dataa(!read_latency_shift_reg_02),
	.datab(!read_latency_shift_reg_03),
	.datac(!read_latency_shift_reg_04),
	.datad(!av_readdata_pre_08),
	.datae(!av_readdata_pre_02),
	.dataf(!av_readdata_pre_03),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[0]~0 .extended_lut = "off";
defparam \src_data[0]~0 .lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam \src_data[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \src_data[0]~3 (
	.dataa(!read_latency_shift_reg_013),
	.datab(!read_latency_shift_reg_015),
	.datac(!av_readdata_pre_06),
	.datad(!av_readdata_pre_014),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[0]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[0]~3 .extended_lut = "off";
defparam \src_data[0]~3 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[0]~3 .shared_arith = "off";

cyclonev_lcell_comb \src_data[0]~4 (
	.dataa(!read_latency_shift_reg_07),
	.datab(!read_latency_shift_reg_08),
	.datac(!av_readdata_pre_015),
	.datad(!av_readdata_pre_016),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[0]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[0]~4 .extended_lut = "off";
defparam \src_data[0]~4 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[0]~4 .shared_arith = "off";

cyclonev_lcell_comb \src_data[0]~5 (
	.dataa(!read_latency_shift_reg_016),
	.datab(!read_latency_shift_reg_09),
	.datac(!av_readdata_pre_05),
	.datad(!av_readdata_pre_013),
	.datae(!\src_data[0]~3_combout ),
	.dataf(!\src_data[0]~4_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[0]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[0]~5 .extended_lut = "off";
defparam \src_data[0]~5 .lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam \src_data[0]~5 .shared_arith = "off";

cyclonev_lcell_comb \src_data[0]~18 (
	.dataa(!read_latency_shift_reg_012),
	.datab(!av_readdata_pre_01),
	.datac(!read_latency_shift_reg_01),
	.datad(!av_readdata_pre_011),
	.datae(!src0_valid),
	.dataf(!av_readdata_pre_07),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[0]~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[0]~18 .extended_lut = "off";
defparam \src_data[0]~18 .lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam \src_data[0]~18 .shared_arith = "off";

cyclonev_lcell_comb \src_data[0]~1 (
	.dataa(!read_latency_shift_reg_05),
	.datab(!read_latency_shift_reg_06),
	.datac(!av_readdata_pre_09),
	.datad(!av_readdata_pre_010),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[0]~1 .extended_lut = "off";
defparam \src_data[0]~1 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \src_data[0]~2 (
	.dataa(!read_latency_shift_reg_010),
	.datab(!read_latency_shift_reg_011),
	.datac(!av_readdata_pre_012),
	.datad(!av_readdata_pre_04),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[0]~2 .extended_lut = "off";
defparam \src_data[0]~2 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[0]~2 .shared_arith = "off";

cyclonev_lcell_comb \src_data[0]~19 (
	.dataa(!\src_data[0]~1_combout ),
	.datab(!\src_data[0]~2_combout ),
	.datac(!read_latency_shift_reg_0),
	.datad(!av_readdata_pre_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[0]~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[0]~19 .extended_lut = "off";
defparam \src_data[0]~19 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \src_data[0]~19 .shared_arith = "off";

cyclonev_lcell_comb \src_data[1]~6 (
	.dataa(!read_latency_shift_reg_013),
	.datab(!read_latency_shift_reg_015),
	.datac(!av_readdata_pre_11),
	.datad(!src_payload),
	.datae(!av_readdata_pre_112),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[1]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[1]~6 .extended_lut = "off";
defparam \src_data[1]~6 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \src_data[1]~6 .shared_arith = "off";

cyclonev_lcell_comb \src_data[1]~7 (
	.dataa(!read_latency_shift_reg_08),
	.datab(!read_latency_shift_reg_01),
	.datac(!av_readdata_pre_113),
	.datad(!av_readdata_pre_114),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[1]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[1]~7 .extended_lut = "off";
defparam \src_data[1]~7 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[1]~7 .shared_arith = "off";

cyclonev_lcell_comb \src_data[1]~20 (
	.dataa(!read_latency_shift_reg_06),
	.datab(!av_readdata_pre_14),
	.datac(!read_latency_shift_reg_07),
	.datad(!av_readdata_pre_110),
	.datae(!read_latency_shift_reg_02),
	.dataf(!av_readdata_pre_111),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[1]~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[1]~20 .extended_lut = "off";
defparam \src_data[1]~20 .lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam \src_data[1]~20 .shared_arith = "off";

cyclonev_lcell_comb \src_data[1]~8 (
	.dataa(!read_latency_shift_reg_03),
	.datab(!read_latency_shift_reg_04),
	.datac(!read_latency_shift_reg_05),
	.datad(!av_readdata_pre_12),
	.datae(!av_readdata_pre_13),
	.dataf(!av_readdata_pre_115),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[1]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[1]~8 .extended_lut = "off";
defparam \src_data[1]~8 .lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam \src_data[1]~8 .shared_arith = "off";

cyclonev_lcell_comb \src_data[1]~21 (
	.dataa(!\src_data[1]~8_combout ),
	.datab(!read_latency_shift_reg_016),
	.datac(!src0_valid),
	.datad(!av_readdata_pre_15),
	.datae(!av_readdata_pre_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[1]~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[1]~21 .extended_lut = "off";
defparam \src_data[1]~21 .lut_mask = 64'hFFFFFFFDFFFFFFFD;
defparam \src_data[1]~21 .shared_arith = "off";

cyclonev_lcell_comb \src_data[2]~9 (
	.dataa(!read_latency_shift_reg_013),
	.datab(!read_latency_shift_reg_015),
	.datac(!src_payload),
	.datad(!av_readdata_pre_21),
	.datae(!av_readdata_pre_28),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[2]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[2]~9 .extended_lut = "off";
defparam \src_data[2]~9 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \src_data[2]~9 .shared_arith = "off";

cyclonev_lcell_comb \src_data[2]~10 (
	.dataa(!read_latency_shift_reg_08),
	.datab(!read_latency_shift_reg_01),
	.datac(!av_readdata_pre_29),
	.datad(!av_readdata_pre_210),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[2]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[2]~10 .extended_lut = "off";
defparam \src_data[2]~10 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[2]~10 .shared_arith = "off";

cyclonev_lcell_comb \src_data[2]~22 (
	.dataa(!read_latency_shift_reg_06),
	.datab(!av_readdata_pre_24),
	.datac(!read_latency_shift_reg_07),
	.datad(!av_readdata_pre_26),
	.datae(!read_latency_shift_reg_02),
	.dataf(!av_readdata_pre_27),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[2]~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[2]~22 .extended_lut = "off";
defparam \src_data[2]~22 .lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam \src_data[2]~22 .shared_arith = "off";

cyclonev_lcell_comb \src_data[2]~11 (
	.dataa(!read_latency_shift_reg_03),
	.datab(!read_latency_shift_reg_04),
	.datac(!read_latency_shift_reg_05),
	.datad(!av_readdata_pre_22),
	.datae(!av_readdata_pre_23),
	.dataf(!av_readdata_pre_212),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[2]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[2]~11 .extended_lut = "off";
defparam \src_data[2]~11 .lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam \src_data[2]~11 .shared_arith = "off";

cyclonev_lcell_comb \src_data[2]~23 (
	.dataa(!\src_data[2]~11_combout ),
	.datab(!read_latency_shift_reg_016),
	.datac(!src0_valid),
	.datad(!av_readdata_pre_25),
	.datae(!av_readdata_pre_2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[2]~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[2]~23 .extended_lut = "off";
defparam \src_data[2]~23 .lut_mask = 64'hFFFFFFFDFFFFFFFD;
defparam \src_data[2]~23 .shared_arith = "off";

cyclonev_lcell_comb \src_data[3]~12 (
	.dataa(!read_latency_shift_reg_07),
	.datab(!src0_valid),
	.datac(!av_readdata_pre_36),
	.datad(!av_readdata_pre_37),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[3]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[3]~12 .extended_lut = "off";
defparam \src_data[3]~12 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[3]~12 .shared_arith = "off";

cyclonev_lcell_comb \src_data[3]~13 (
	.dataa(!read_latency_shift_reg_04),
	.datab(!read_latency_shift_reg_05),
	.datac(!av_readdata_pre_3),
	.datad(!av_readdata_pre_38),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[3]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[3]~13 .extended_lut = "off";
defparam \src_data[3]~13 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[3]~13 .shared_arith = "off";

cyclonev_lcell_comb \src_data[3]~14 (
	.dataa(!read_latency_shift_reg_013),
	.datab(!read_latency_shift_reg_015),
	.datac(!av_readdata_pre_33),
	.datad(!av_readdata_pre_39),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[3]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[3]~14 .extended_lut = "off";
defparam \src_data[3]~14 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[3]~14 .shared_arith = "off";

cyclonev_lcell_comb \src_data[3]~15 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!read_latency_shift_reg_02),
	.datac(!av_readdata_pre_310),
	.datad(!av_readdata_pre_311),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[3]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[3]~15 .extended_lut = "off";
defparam \src_data[3]~15 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[3]~15 .shared_arith = "off";

cyclonev_lcell_comb \src_data[3]~16 (
	.dataa(!read_latency_shift_reg_016),
	.datab(!read_latency_shift_reg_03),
	.datac(!av_readdata_pre_31),
	.datad(!av_readdata_pre_32),
	.datae(!\src_data[3]~14_combout ),
	.dataf(!\src_data[3]~15_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[3]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[3]~16 .extended_lut = "off";
defparam \src_data[3]~16 .lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam \src_data[3]~16 .shared_arith = "off";

cyclonev_lcell_comb \src_data[3]~17 (
	.dataa(!read_latency_shift_reg_06),
	.datab(!av_readdata_pre_35),
	.datac(!\src_data[3]~12_combout ),
	.datad(!\src_data[3]~13_combout ),
	.datae(!\src_data[3]~16_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[3]~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[3]~17 .extended_lut = "off";
defparam \src_data[3]~17 .lut_mask = 64'hFFFEFFFFFFFEFFFF;
defparam \src_data[3]~17 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~1 (
	.dataa(!read_latency_shift_reg_08),
	.datab(!read_latency_shift_reg_01),
	.datac(!read_latency_shift_reg_02),
	.datad(!av_readdata_pre_47),
	.datae(!av_readdata_pre_48),
	.dataf(!av_readdata_pre_49),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~1 .extended_lut = "off";
defparam \src_payload~1 .lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam \src_payload~1 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~2 (
	.dataa(!read_latency_shift_reg_03),
	.datab(!read_latency_shift_reg_04),
	.datac(!av_readdata_pre_42),
	.datad(!av_readdata_pre_43),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~2 .extended_lut = "off";
defparam \src_payload~2 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_payload~2 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~52 (
	.dataa(!read_latency_shift_reg_07),
	.datab(!av_readdata_pre_46),
	.datac(!read_latency_shift_reg_015),
	.datad(!av_readdata_pre_44),
	.datae(!src0_valid),
	.dataf(!av_readdata_pre_45),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~52_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~52 .extended_lut = "off";
defparam \src_payload~52 .lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam \src_payload~52 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~53 (
	.dataa(!read_latency_shift_reg_013),
	.datab(!src_payload),
	.datac(!av_readdata_pre_4),
	.datad(!read_latency_shift_reg_016),
	.datae(!av_readdata_pre_41),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~53_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~53 .extended_lut = "off";
defparam \src_payload~53 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \src_payload~53 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~4 (
	.dataa(!read_latency_shift_reg_013),
	.datab(!read_latency_shift_reg_015),
	.datac(!av_readdata_pre_53),
	.datad(!av_readdata_pre_57),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~4 .extended_lut = "off";
defparam \src_payload~4 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_payload~4 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~5 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!read_latency_shift_reg_02),
	.datac(!av_readdata_pre_58),
	.datad(!av_readdata_pre_59),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~5 .extended_lut = "off";
defparam \src_payload~5 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_payload~5 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~6 (
	.dataa(!read_latency_shift_reg_016),
	.datab(!read_latency_shift_reg_03),
	.datac(!av_readdata_pre_51),
	.datad(!av_readdata_pre_52),
	.datae(!\src_payload~4_combout ),
	.dataf(!\src_payload~5_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~6 .extended_lut = "off";
defparam \src_payload~6 .lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam \src_payload~6 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~54 (
	.dataa(!read_latency_shift_reg_04),
	.datab(!av_readdata_pre_5),
	.datac(!read_latency_shift_reg_08),
	.datad(!av_readdata_pre_56),
	.datae(!src0_valid),
	.dataf(!av_readdata_pre_54),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~54_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~54 .extended_lut = "off";
defparam \src_payload~54 .lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam \src_payload~54 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~8 (
	.dataa(!read_latency_shift_reg_013),
	.datab(!read_latency_shift_reg_015),
	.datac(!src_payload),
	.datad(!av_readdata_pre_61),
	.datae(!av_readdata_pre_65),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~8 .extended_lut = "off";
defparam \src_payload~8 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \src_payload~8 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~9 (
	.dataa(!read_latency_shift_reg_016),
	.datab(!src0_valid),
	.datac(!av_readdata_pre_66),
	.datad(!av_readdata_pre_62),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~9 .extended_lut = "off";
defparam \src_payload~9 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_payload~9 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~10 (
	.dataa(!read_latency_shift_reg_08),
	.datab(!read_latency_shift_reg_03),
	.datac(!av_readdata_pre_67),
	.datad(!av_readdata_pre_63),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~10 .extended_lut = "off";
defparam \src_payload~10 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_payload~10 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~11 (
	.dataa(!read_latency_shift_reg_04),
	.datab(!av_readdata_pre_6),
	.datac(!\src_payload~8_combout ),
	.datad(!\src_payload~9_combout ),
	.datae(!\src_payload~10_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~11 .extended_lut = "off";
defparam \src_payload~11 .lut_mask = 64'hFFFFFFEFFFFFFFEF;
defparam \src_payload~11 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~13 (
	.dataa(!read_latency_shift_reg_013),
	.datab(!read_latency_shift_reg_015),
	.datac(!src_payload),
	.datad(!av_readdata_pre_7),
	.datae(!av_readdata_pre_72),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~13 .extended_lut = "off";
defparam \src_payload~13 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \src_payload~13 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~14 (
	.dataa(!read_latency_shift_reg_016),
	.datab(!src0_valid),
	.datac(!av_readdata_pre_73),
	.datad(!av_readdata_pre_71),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~14 .extended_lut = "off";
defparam \src_payload~14 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_payload~14 .shared_arith = "off";

endmodule

module first_nios2_system_first_nios2_system_mm_interconnect_0_rsp_mux_001 (
	q_a_0,
	q_a_1,
	q_a_2,
	q_a_3,
	q_a_4,
	q_a_5,
	q_a_6,
	q_a_7,
	q_a_22,
	q_a_23,
	q_a_24,
	q_a_25,
	q_a_31,
	q_a_21,
	q_a_11,
	q_a_28,
	q_a_10,
	q_a_27,
	q_a_8,
	q_a_9,
	q_a_26,
	q_a_20,
	q_a_19,
	q_a_17,
	q_a_30,
	q_a_18,
	q_a_16,
	q_a_15,
	q_a_12,
	q_a_13,
	q_a_14,
	q_a_29,
	src1_valid,
	src1_valid1,
	av_readdata_pre_0,
	av_readdata_pre_1,
	av_readdata_pre_2,
	av_readdata_pre_3,
	av_readdata_pre_4,
	av_readdata_pre_5,
	av_readdata_pre_6,
	av_readdata_pre_7,
	av_readdata_pre_22,
	av_readdata_pre_23,
	av_readdata_pre_24,
	av_readdata_pre_25,
	av_readdata_pre_31,
	av_readdata_pre_21,
	av_readdata_pre_11,
	av_readdata_pre_28,
	av_readdata_pre_10,
	av_readdata_pre_27,
	av_readdata_pre_8,
	av_readdata_pre_9,
	av_readdata_pre_26,
	av_readdata_pre_20,
	av_readdata_pre_19,
	av_readdata_pre_17,
	av_readdata_pre_30,
	av_readdata_pre_18,
	av_readdata_pre_16,
	av_readdata_pre_15,
	av_readdata_pre_12,
	av_readdata_pre_13,
	av_readdata_pre_14,
	av_readdata_pre_29,
	WideOr11,
	src_data_26,
	src_data_25,
	src_data_24,
	src_data_23,
	src_data_22,
	src_data_1,
	src_data_0,
	src_data_2,
	src_data_3,
	src_data_4,
	src_data_5,
	src_data_28,
	src_data_31,
	src_data_27,
	src_data_29,
	src_data_30,
	src_data_11,
	src_data_12,
	src_data_13,
	src_data_14,
	src_data_15,
	src_data_16,
	src_data_9,
	src_data_21,
	src_data_6,
	src_data_8,
	src_data_17,
	src_data_18,
	src_data_10,
	src_data_7,
	src_data_20,
	src_data_19)/* synthesis synthesis_greybox=1 */;
input 	q_a_0;
input 	q_a_1;
input 	q_a_2;
input 	q_a_3;
input 	q_a_4;
input 	q_a_5;
input 	q_a_6;
input 	q_a_7;
input 	q_a_22;
input 	q_a_23;
input 	q_a_24;
input 	q_a_25;
input 	q_a_31;
input 	q_a_21;
input 	q_a_11;
input 	q_a_28;
input 	q_a_10;
input 	q_a_27;
input 	q_a_8;
input 	q_a_9;
input 	q_a_26;
input 	q_a_20;
input 	q_a_19;
input 	q_a_17;
input 	q_a_30;
input 	q_a_18;
input 	q_a_16;
input 	q_a_15;
input 	q_a_12;
input 	q_a_13;
input 	q_a_14;
input 	q_a_29;
input 	src1_valid;
input 	src1_valid1;
input 	av_readdata_pre_0;
input 	av_readdata_pre_1;
input 	av_readdata_pre_2;
input 	av_readdata_pre_3;
input 	av_readdata_pre_4;
input 	av_readdata_pre_5;
input 	av_readdata_pre_6;
input 	av_readdata_pre_7;
input 	av_readdata_pre_22;
input 	av_readdata_pre_23;
input 	av_readdata_pre_24;
input 	av_readdata_pre_25;
input 	av_readdata_pre_31;
input 	av_readdata_pre_21;
input 	av_readdata_pre_11;
input 	av_readdata_pre_28;
input 	av_readdata_pre_10;
input 	av_readdata_pre_27;
input 	av_readdata_pre_8;
input 	av_readdata_pre_9;
input 	av_readdata_pre_26;
input 	av_readdata_pre_20;
input 	av_readdata_pre_19;
input 	av_readdata_pre_17;
input 	av_readdata_pre_30;
input 	av_readdata_pre_18;
input 	av_readdata_pre_16;
input 	av_readdata_pre_15;
input 	av_readdata_pre_12;
input 	av_readdata_pre_13;
input 	av_readdata_pre_14;
input 	av_readdata_pre_29;
output 	WideOr11;
output 	src_data_26;
output 	src_data_25;
output 	src_data_24;
output 	src_data_23;
output 	src_data_22;
output 	src_data_1;
output 	src_data_0;
output 	src_data_2;
output 	src_data_3;
output 	src_data_4;
output 	src_data_5;
output 	src_data_28;
output 	src_data_31;
output 	src_data_27;
output 	src_data_29;
output 	src_data_30;
output 	src_data_11;
output 	src_data_12;
output 	src_data_13;
output 	src_data_14;
output 	src_data_15;
output 	src_data_16;
output 	src_data_9;
output 	src_data_21;
output 	src_data_6;
output 	src_data_8;
output 	src_data_17;
output 	src_data_18;
output 	src_data_10;
output 	src_data_7;
output 	src_data_20;
output 	src_data_19;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb WideOr1(
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr11),
	.sumout(),
	.cout(),
	.shareout());
defparam WideOr1.extended_lut = "off";
defparam WideOr1.lut_mask = 64'h7777777777777777;
defparam WideOr1.shared_arith = "off";

cyclonev_lcell_comb \src_data[26] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_26),
	.datad(!q_a_26),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_26),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[26] .extended_lut = "off";
defparam \src_data[26] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[26] .shared_arith = "off";

cyclonev_lcell_comb \src_data[25] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_25),
	.datad(!q_a_25),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_25),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[25] .extended_lut = "off";
defparam \src_data[25] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[25] .shared_arith = "off";

cyclonev_lcell_comb \src_data[24] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_24),
	.datad(!q_a_24),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_24),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[24] .extended_lut = "off";
defparam \src_data[24] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[24] .shared_arith = "off";

cyclonev_lcell_comb \src_data[23] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_23),
	.datad(!q_a_23),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_23),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[23] .extended_lut = "off";
defparam \src_data[23] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[23] .shared_arith = "off";

cyclonev_lcell_comb \src_data[22] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_22),
	.datad(!q_a_22),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_22),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[22] .extended_lut = "off";
defparam \src_data[22] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[22] .shared_arith = "off";

cyclonev_lcell_comb \src_data[1] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_1),
	.datad(!q_a_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[1] .extended_lut = "off";
defparam \src_data[1] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[1] .shared_arith = "off";

cyclonev_lcell_comb \src_data[0] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_0),
	.datad(!q_a_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[0] .extended_lut = "off";
defparam \src_data[0] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[0] .shared_arith = "off";

cyclonev_lcell_comb \src_data[2] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_2),
	.datad(!q_a_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_2),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[2] .extended_lut = "off";
defparam \src_data[2] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[2] .shared_arith = "off";

cyclonev_lcell_comb \src_data[3] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_3),
	.datad(!q_a_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_3),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[3] .extended_lut = "off";
defparam \src_data[3] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[3] .shared_arith = "off";

cyclonev_lcell_comb \src_data[4] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_4),
	.datad(!q_a_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_4),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[4] .extended_lut = "off";
defparam \src_data[4] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[4] .shared_arith = "off";

cyclonev_lcell_comb \src_data[5] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_5),
	.datad(!q_a_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_5),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[5] .extended_lut = "off";
defparam \src_data[5] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[5] .shared_arith = "off";

cyclonev_lcell_comb \src_data[28] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_28),
	.datad(!q_a_28),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_28),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[28] .extended_lut = "off";
defparam \src_data[28] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[28] .shared_arith = "off";

cyclonev_lcell_comb \src_data[31] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_31),
	.datad(!q_a_31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_31),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[31] .extended_lut = "off";
defparam \src_data[31] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[31] .shared_arith = "off";

cyclonev_lcell_comb \src_data[27] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_27),
	.datad(!q_a_27),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_27),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[27] .extended_lut = "off";
defparam \src_data[27] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[27] .shared_arith = "off";

cyclonev_lcell_comb \src_data[29] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_29),
	.datad(!q_a_29),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_29),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[29] .extended_lut = "off";
defparam \src_data[29] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[29] .shared_arith = "off";

cyclonev_lcell_comb \src_data[30] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_30),
	.datad(!q_a_30),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_30),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[30] .extended_lut = "off";
defparam \src_data[30] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[30] .shared_arith = "off";

cyclonev_lcell_comb \src_data[11] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_11),
	.datad(!q_a_11),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_11),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[11] .extended_lut = "off";
defparam \src_data[11] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[11] .shared_arith = "off";

cyclonev_lcell_comb \src_data[12] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_12),
	.datad(!q_a_12),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_12),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[12] .extended_lut = "off";
defparam \src_data[12] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[12] .shared_arith = "off";

cyclonev_lcell_comb \src_data[13] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_13),
	.datad(!q_a_13),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_13),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[13] .extended_lut = "off";
defparam \src_data[13] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[13] .shared_arith = "off";

cyclonev_lcell_comb \src_data[14] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_14),
	.datad(!q_a_14),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_14),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[14] .extended_lut = "off";
defparam \src_data[14] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[14] .shared_arith = "off";

cyclonev_lcell_comb \src_data[15] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_15),
	.datad(!q_a_15),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_15),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[15] .extended_lut = "off";
defparam \src_data[15] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[15] .shared_arith = "off";

cyclonev_lcell_comb \src_data[16] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_16),
	.datad(!q_a_16),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_16),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[16] .extended_lut = "off";
defparam \src_data[16] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[16] .shared_arith = "off";

cyclonev_lcell_comb \src_data[9] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_9),
	.datad(!q_a_9),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_9),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[9] .extended_lut = "off";
defparam \src_data[9] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[9] .shared_arith = "off";

cyclonev_lcell_comb \src_data[21] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_21),
	.datad(!q_a_21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_21),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[21] .extended_lut = "off";
defparam \src_data[21] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[21] .shared_arith = "off";

cyclonev_lcell_comb \src_data[6] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_6),
	.datad(!q_a_6),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_6),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[6] .extended_lut = "off";
defparam \src_data[6] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[6] .shared_arith = "off";

cyclonev_lcell_comb \src_data[8] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_8),
	.datad(!q_a_8),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_8),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[8] .extended_lut = "off";
defparam \src_data[8] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[8] .shared_arith = "off";

cyclonev_lcell_comb \src_data[17] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_17),
	.datad(!q_a_17),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_17),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[17] .extended_lut = "off";
defparam \src_data[17] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[17] .shared_arith = "off";

cyclonev_lcell_comb \src_data[18] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_18),
	.datad(!q_a_18),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_18),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[18] .extended_lut = "off";
defparam \src_data[18] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[18] .shared_arith = "off";

cyclonev_lcell_comb \src_data[10] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_10),
	.datad(!q_a_10),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_10),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[10] .extended_lut = "off";
defparam \src_data[10] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[10] .shared_arith = "off";

cyclonev_lcell_comb \src_data[7] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_7),
	.datad(!q_a_7),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_7),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[7] .extended_lut = "off";
defparam \src_data[7] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[7] .shared_arith = "off";

cyclonev_lcell_comb \src_data[20] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_20),
	.datad(!q_a_20),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_20),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[20] .extended_lut = "off";
defparam \src_data[20] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[20] .shared_arith = "off";

cyclonev_lcell_comb \src_data[19] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_19),
	.datad(!q_a_19),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_19),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[19] .extended_lut = "off";
defparam \src_data[19] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[19] .shared_arith = "off";

endmodule

module first_nios2_system_first_nios2_system_onchip_mem (
	q_a_0,
	q_a_1,
	q_a_2,
	q_a_3,
	q_a_4,
	q_a_5,
	q_a_6,
	q_a_7,
	q_a_22,
	q_a_23,
	q_a_24,
	q_a_25,
	q_a_31,
	q_a_21,
	q_a_11,
	q_a_28,
	q_a_10,
	q_a_27,
	q_a_8,
	q_a_9,
	q_a_26,
	q_a_20,
	q_a_19,
	q_a_17,
	q_a_30,
	q_a_18,
	q_a_16,
	q_a_15,
	q_a_12,
	q_a_13,
	q_a_14,
	q_a_29,
	d_write,
	mem_used_1,
	saved_grant_0,
	WideOr1,
	r_early_rst,
	src_payload,
	src_data_38,
	src_data_39,
	src_data_40,
	src_data_41,
	src_data_42,
	src_data_43,
	src_data_44,
	src_data_45,
	src_data_46,
	src_data_47,
	src_data_48,
	src_data_49,
	src_data_50,
	src_data_32,
	src_payload1,
	src_payload2,
	src_payload3,
	src_payload4,
	src_payload5,
	src_payload6,
	src_payload7,
	src_payload8,
	src_data_34,
	src_payload9,
	src_payload10,
	src_data_35,
	src_payload11,
	src_payload12,
	src_payload13,
	src_payload14,
	src_data_33,
	src_payload15,
	src_payload16,
	src_payload17,
	src_payload18,
	src_payload19,
	src_payload20,
	src_payload21,
	src_payload22,
	src_payload23,
	src_payload24,
	src_payload25,
	src_payload26,
	src_payload27,
	src_payload28,
	src_payload29,
	src_payload30,
	src_payload31,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	q_a_0;
output 	q_a_1;
output 	q_a_2;
output 	q_a_3;
output 	q_a_4;
output 	q_a_5;
output 	q_a_6;
output 	q_a_7;
output 	q_a_22;
output 	q_a_23;
output 	q_a_24;
output 	q_a_25;
output 	q_a_31;
output 	q_a_21;
output 	q_a_11;
output 	q_a_28;
output 	q_a_10;
output 	q_a_27;
output 	q_a_8;
output 	q_a_9;
output 	q_a_26;
output 	q_a_20;
output 	q_a_19;
output 	q_a_17;
output 	q_a_30;
output 	q_a_18;
output 	q_a_16;
output 	q_a_15;
output 	q_a_12;
output 	q_a_13;
output 	q_a_14;
output 	q_a_29;
input 	d_write;
input 	mem_used_1;
input 	saved_grant_0;
input 	WideOr1;
input 	r_early_rst;
input 	src_payload;
input 	src_data_38;
input 	src_data_39;
input 	src_data_40;
input 	src_data_41;
input 	src_data_42;
input 	src_data_43;
input 	src_data_44;
input 	src_data_45;
input 	src_data_46;
input 	src_data_47;
input 	src_data_48;
input 	src_data_49;
input 	src_data_50;
input 	src_data_32;
input 	src_payload1;
input 	src_payload2;
input 	src_payload3;
input 	src_payload4;
input 	src_payload5;
input 	src_payload6;
input 	src_payload7;
input 	src_payload8;
input 	src_data_34;
input 	src_payload9;
input 	src_payload10;
input 	src_data_35;
input 	src_payload11;
input 	src_payload12;
input 	src_payload13;
input 	src_payload14;
input 	src_data_33;
input 	src_payload15;
input 	src_payload16;
input 	src_payload17;
input 	src_payload18;
input 	src_payload19;
input 	src_payload20;
input 	src_payload21;
input 	src_payload22;
input 	src_payload23;
input 	src_payload24;
input 	src_payload25;
input 	src_payload26;
input 	src_payload27;
input 	src_payload28;
input 	src_payload29;
input 	src_payload30;
input 	src_payload31;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wren~0_combout ;


first_nios2_system_altsyncram_7 the_altsyncram(
	.q_a({q_a_31,q_a_30,q_a_29,q_a_28,q_a_27,q_a_26,q_a_25,q_a_24,q_a_23,q_a_22,q_a_21,q_a_20,q_a_19,q_a_18,q_a_17,q_a_16,q_a_15,q_a_14,q_a_13,q_a_12,q_a_11,q_a_10,q_a_9,q_a_8,q_a_7,q_a_6,q_a_5,q_a_4,q_a_3,q_a_2,q_a_1,q_a_0}),
	.clocken0(r_early_rst),
	.wren_a(\wren~0_combout ),
	.data_a({src_payload12,src_payload24,src_payload31,src_payload15,src_payload17,src_payload20,src_payload11,src_payload10,src_payload9,src_payload8,src_payload13,src_payload21,src_payload22,src_payload25,src_payload23,src_payload26,src_payload27,src_payload30,src_payload29,
src_payload28,src_payload14,src_payload16,src_payload19,src_payload18,src_payload7,src_payload6,src_payload5,src_payload4,src_payload3,src_payload2,src_payload1,src_payload}),
	.address_a({src_data_50,src_data_49,src_data_48,src_data_47,src_data_46,src_data_45,src_data_44,src_data_43,src_data_42,src_data_41,src_data_40,src_data_39,src_data_38}),
	.byteena_a({src_data_35,src_data_34,src_data_33,src_data_32}),
	.clock0(clk_clk));

cyclonev_lcell_comb \wren~0 (
	.dataa(!d_write),
	.datab(!mem_used_1),
	.datac(!saved_grant_0),
	.datad(!WideOr1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wren~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wren~0 .extended_lut = "off";
defparam \wren~0 .lut_mask = 64'hFBFFFBFFFBFFFBFF;
defparam \wren~0 .shared_arith = "off";

endmodule

module first_nios2_system_altsyncram_7 (
	q_a,
	clocken0,
	wren_a,
	data_a,
	address_a,
	byteena_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_a;
input 	clocken0;
input 	wren_a;
input 	[31:0] data_a;
input 	[12:0] address_a;
input 	[3:0] byteena_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



first_nios2_system_altsyncram_mun1 auto_generated(
	.q_a({q_a[31],q_a[30],q_a[29],q_a[28],q_a[27],q_a[26],q_a[25],q_a[24],q_a[23],q_a[22],q_a[21],q_a[20],q_a[19],q_a[18],q_a[17],q_a[16],q_a[15],q_a[14],q_a[13],q_a[12],q_a[11],q_a[10],q_a[9],q_a[8],q_a[7],q_a[6],q_a[5],q_a[4],q_a[3],q_a[2],q_a[1],q_a[0]}),
	.clocken0(clocken0),
	.wren_a(wren_a),
	.data_a({data_a[31],data_a[30],data_a[29],data_a[28],data_a[27],data_a[26],data_a[25],data_a[24],data_a[23],data_a[22],data_a[21],data_a[20],data_a[19],data_a[18],data_a[17],data_a[16],data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.address_a({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.byteena_a({byteena_a[3],byteena_a[2],byteena_a[1],byteena_a[0]}),
	.clock0(clock0));

endmodule

module first_nios2_system_altsyncram_mun1 (
	q_a,
	clocken0,
	wren_a,
	data_a,
	address_a,
	byteena_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_a;
input 	clocken0;
input 	wren_a;
input 	[31:0] data_a;
input 	[12:0] address_a;
input 	[3:0] byteena_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTADATAOUT_bus;
wire [143:0] ram_block1a1_PORTADATAOUT_bus;
wire [143:0] ram_block1a2_PORTADATAOUT_bus;
wire [143:0] ram_block1a3_PORTADATAOUT_bus;
wire [143:0] ram_block1a4_PORTADATAOUT_bus;
wire [143:0] ram_block1a5_PORTADATAOUT_bus;
wire [143:0] ram_block1a6_PORTADATAOUT_bus;
wire [143:0] ram_block1a7_PORTADATAOUT_bus;
wire [143:0] ram_block1a22_PORTADATAOUT_bus;
wire [143:0] ram_block1a23_PORTADATAOUT_bus;
wire [143:0] ram_block1a24_PORTADATAOUT_bus;
wire [143:0] ram_block1a25_PORTADATAOUT_bus;
wire [143:0] ram_block1a31_PORTADATAOUT_bus;
wire [143:0] ram_block1a21_PORTADATAOUT_bus;
wire [143:0] ram_block1a11_PORTADATAOUT_bus;
wire [143:0] ram_block1a28_PORTADATAOUT_bus;
wire [143:0] ram_block1a10_PORTADATAOUT_bus;
wire [143:0] ram_block1a27_PORTADATAOUT_bus;
wire [143:0] ram_block1a8_PORTADATAOUT_bus;
wire [143:0] ram_block1a9_PORTADATAOUT_bus;
wire [143:0] ram_block1a26_PORTADATAOUT_bus;
wire [143:0] ram_block1a20_PORTADATAOUT_bus;
wire [143:0] ram_block1a19_PORTADATAOUT_bus;
wire [143:0] ram_block1a17_PORTADATAOUT_bus;
wire [143:0] ram_block1a30_PORTADATAOUT_bus;
wire [143:0] ram_block1a18_PORTADATAOUT_bus;
wire [143:0] ram_block1a16_PORTADATAOUT_bus;
wire [143:0] ram_block1a15_PORTADATAOUT_bus;
wire [143:0] ram_block1a12_PORTADATAOUT_bus;
wire [143:0] ram_block1a13_PORTADATAOUT_bus;
wire [143:0] ram_block1a14_PORTADATAOUT_bus;
wire [143:0] ram_block1a29_PORTADATAOUT_bus;

assign q_a[0] = ram_block1a0_PORTADATAOUT_bus[0];

assign q_a[1] = ram_block1a1_PORTADATAOUT_bus[0];

assign q_a[2] = ram_block1a2_PORTADATAOUT_bus[0];

assign q_a[3] = ram_block1a3_PORTADATAOUT_bus[0];

assign q_a[4] = ram_block1a4_PORTADATAOUT_bus[0];

assign q_a[5] = ram_block1a5_PORTADATAOUT_bus[0];

assign q_a[6] = ram_block1a6_PORTADATAOUT_bus[0];

assign q_a[7] = ram_block1a7_PORTADATAOUT_bus[0];

assign q_a[22] = ram_block1a22_PORTADATAOUT_bus[0];

assign q_a[23] = ram_block1a23_PORTADATAOUT_bus[0];

assign q_a[24] = ram_block1a24_PORTADATAOUT_bus[0];

assign q_a[25] = ram_block1a25_PORTADATAOUT_bus[0];

assign q_a[31] = ram_block1a31_PORTADATAOUT_bus[0];

assign q_a[21] = ram_block1a21_PORTADATAOUT_bus[0];

assign q_a[11] = ram_block1a11_PORTADATAOUT_bus[0];

assign q_a[28] = ram_block1a28_PORTADATAOUT_bus[0];

assign q_a[10] = ram_block1a10_PORTADATAOUT_bus[0];

assign q_a[27] = ram_block1a27_PORTADATAOUT_bus[0];

assign q_a[8] = ram_block1a8_PORTADATAOUT_bus[0];

assign q_a[9] = ram_block1a9_PORTADATAOUT_bus[0];

assign q_a[26] = ram_block1a26_PORTADATAOUT_bus[0];

assign q_a[20] = ram_block1a20_PORTADATAOUT_bus[0];

assign q_a[19] = ram_block1a19_PORTADATAOUT_bus[0];

assign q_a[17] = ram_block1a17_PORTADATAOUT_bus[0];

assign q_a[30] = ram_block1a30_PORTADATAOUT_bus[0];

assign q_a[18] = ram_block1a18_PORTADATAOUT_bus[0];

assign q_a[16] = ram_block1a16_PORTADATAOUT_bus[0];

assign q_a[15] = ram_block1a15_PORTADATAOUT_bus[0];

assign q_a[12] = ram_block1a12_PORTADATAOUT_bus[0];

assign q_a[13] = ram_block1a13_PORTADATAOUT_bus[0];

assign q_a[14] = ram_block1a14_PORTADATAOUT_bus[0];

assign q_a[29] = ram_block1a29_PORTADATAOUT_bus[0];

cyclonev_ram_block ram_block1a0(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a0_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.init_file = "first_nios2_system_onchip_mem.hex";
defparam ram_block1a0.init_file_layout = "port_a";
defparam ram_block1a0.logical_ram_name = "first_nios2_system_onchip_mem:onchip_mem|altsyncram:the_altsyncram|altsyncram_mun1:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.operation_mode = "single_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 13;
defparam ram_block1a0.port_a_byte_enable_mask_width = 1;
defparam ram_block1a0.port_a_byte_size = 1;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 5119;
defparam ram_block1a0.port_a_logical_ram_depth = 5120;
defparam ram_block1a0.port_a_logical_ram_width = 32;
defparam ram_block1a0.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a0.ram_block_type = "auto";
defparam ram_block1a0.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a0.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a0.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a1(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a1_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.init_file = "first_nios2_system_onchip_mem.hex";
defparam ram_block1a1.init_file_layout = "port_a";
defparam ram_block1a1.logical_ram_name = "first_nios2_system_onchip_mem:onchip_mem|altsyncram:the_altsyncram|altsyncram_mun1:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.operation_mode = "single_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 13;
defparam ram_block1a1.port_a_byte_enable_mask_width = 1;
defparam ram_block1a1.port_a_byte_size = 1;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 5119;
defparam ram_block1a1.port_a_logical_ram_depth = 5120;
defparam ram_block1a1.port_a_logical_ram_width = 32;
defparam ram_block1a1.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a1.ram_block_type = "auto";
defparam ram_block1a1.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a1.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a1.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a2(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a2_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.init_file = "first_nios2_system_onchip_mem.hex";
defparam ram_block1a2.init_file_layout = "port_a";
defparam ram_block1a2.logical_ram_name = "first_nios2_system_onchip_mem:onchip_mem|altsyncram:the_altsyncram|altsyncram_mun1:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.operation_mode = "single_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 13;
defparam ram_block1a2.port_a_byte_enable_mask_width = 1;
defparam ram_block1a2.port_a_byte_size = 1;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 5119;
defparam ram_block1a2.port_a_logical_ram_depth = 5120;
defparam ram_block1a2.port_a_logical_ram_width = 32;
defparam ram_block1a2.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a2.ram_block_type = "auto";
defparam ram_block1a2.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a2.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a2.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a3(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a3_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.init_file = "first_nios2_system_onchip_mem.hex";
defparam ram_block1a3.init_file_layout = "port_a";
defparam ram_block1a3.logical_ram_name = "first_nios2_system_onchip_mem:onchip_mem|altsyncram:the_altsyncram|altsyncram_mun1:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.operation_mode = "single_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 13;
defparam ram_block1a3.port_a_byte_enable_mask_width = 1;
defparam ram_block1a3.port_a_byte_size = 1;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 5119;
defparam ram_block1a3.port_a_logical_ram_depth = 5120;
defparam ram_block1a3.port_a_logical_ram_width = 32;
defparam ram_block1a3.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a3.ram_block_type = "auto";
defparam ram_block1a3.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a3.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a3.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a4(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a4_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.init_file = "first_nios2_system_onchip_mem.hex";
defparam ram_block1a4.init_file_layout = "port_a";
defparam ram_block1a4.logical_ram_name = "first_nios2_system_onchip_mem:onchip_mem|altsyncram:the_altsyncram|altsyncram_mun1:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.operation_mode = "single_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 13;
defparam ram_block1a4.port_a_byte_enable_mask_width = 1;
defparam ram_block1a4.port_a_byte_size = 1;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 5119;
defparam ram_block1a4.port_a_logical_ram_depth = 5120;
defparam ram_block1a4.port_a_logical_ram_width = 32;
defparam ram_block1a4.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a4.ram_block_type = "auto";
defparam ram_block1a4.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a4.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a4.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a5(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a5_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.init_file = "first_nios2_system_onchip_mem.hex";
defparam ram_block1a5.init_file_layout = "port_a";
defparam ram_block1a5.logical_ram_name = "first_nios2_system_onchip_mem:onchip_mem|altsyncram:the_altsyncram|altsyncram_mun1:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.operation_mode = "single_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 13;
defparam ram_block1a5.port_a_byte_enable_mask_width = 1;
defparam ram_block1a5.port_a_byte_size = 1;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 5119;
defparam ram_block1a5.port_a_logical_ram_depth = 5120;
defparam ram_block1a5.port_a_logical_ram_width = 32;
defparam ram_block1a5.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a5.ram_block_type = "auto";
defparam ram_block1a5.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a5.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a5.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a6(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a6_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.init_file = "first_nios2_system_onchip_mem.hex";
defparam ram_block1a6.init_file_layout = "port_a";
defparam ram_block1a6.logical_ram_name = "first_nios2_system_onchip_mem:onchip_mem|altsyncram:the_altsyncram|altsyncram_mun1:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.operation_mode = "single_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 13;
defparam ram_block1a6.port_a_byte_enable_mask_width = 1;
defparam ram_block1a6.port_a_byte_size = 1;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 5119;
defparam ram_block1a6.port_a_logical_ram_depth = 5120;
defparam ram_block1a6.port_a_logical_ram_width = 32;
defparam ram_block1a6.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a6.ram_block_type = "auto";
defparam ram_block1a6.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a6.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a6.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a7(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a7_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.init_file = "first_nios2_system_onchip_mem.hex";
defparam ram_block1a7.init_file_layout = "port_a";
defparam ram_block1a7.logical_ram_name = "first_nios2_system_onchip_mem:onchip_mem|altsyncram:the_altsyncram|altsyncram_mun1:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.operation_mode = "single_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 13;
defparam ram_block1a7.port_a_byte_enable_mask_width = 1;
defparam ram_block1a7.port_a_byte_size = 1;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 5119;
defparam ram_block1a7.port_a_logical_ram_depth = 5120;
defparam ram_block1a7.port_a_logical_ram_width = 32;
defparam ram_block1a7.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a7.ram_block_type = "auto";
defparam ram_block1a7.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a7.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a7.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a22(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[22]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a22_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a22.clk0_core_clock_enable = "ena0";
defparam ram_block1a22.clk0_input_clock_enable = "ena0";
defparam ram_block1a22.data_interleave_offset_in_bits = 1;
defparam ram_block1a22.data_interleave_width_in_bits = 1;
defparam ram_block1a22.init_file = "first_nios2_system_onchip_mem.hex";
defparam ram_block1a22.init_file_layout = "port_a";
defparam ram_block1a22.logical_ram_name = "first_nios2_system_onchip_mem:onchip_mem|altsyncram:the_altsyncram|altsyncram_mun1:auto_generated|ALTSYNCRAM";
defparam ram_block1a22.operation_mode = "single_port";
defparam ram_block1a22.port_a_address_clear = "none";
defparam ram_block1a22.port_a_address_width = 13;
defparam ram_block1a22.port_a_byte_enable_mask_width = 1;
defparam ram_block1a22.port_a_byte_size = 1;
defparam ram_block1a22.port_a_data_out_clear = "none";
defparam ram_block1a22.port_a_data_out_clock = "none";
defparam ram_block1a22.port_a_data_width = 1;
defparam ram_block1a22.port_a_first_address = 0;
defparam ram_block1a22.port_a_first_bit_number = 22;
defparam ram_block1a22.port_a_last_address = 5119;
defparam ram_block1a22.port_a_logical_ram_depth = 5120;
defparam ram_block1a22.port_a_logical_ram_width = 32;
defparam ram_block1a22.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a22.ram_block_type = "auto";
defparam ram_block1a22.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a22.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a22.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a23(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[23]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a23_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a23.clk0_core_clock_enable = "ena0";
defparam ram_block1a23.clk0_input_clock_enable = "ena0";
defparam ram_block1a23.data_interleave_offset_in_bits = 1;
defparam ram_block1a23.data_interleave_width_in_bits = 1;
defparam ram_block1a23.init_file = "first_nios2_system_onchip_mem.hex";
defparam ram_block1a23.init_file_layout = "port_a";
defparam ram_block1a23.logical_ram_name = "first_nios2_system_onchip_mem:onchip_mem|altsyncram:the_altsyncram|altsyncram_mun1:auto_generated|ALTSYNCRAM";
defparam ram_block1a23.operation_mode = "single_port";
defparam ram_block1a23.port_a_address_clear = "none";
defparam ram_block1a23.port_a_address_width = 13;
defparam ram_block1a23.port_a_byte_enable_mask_width = 1;
defparam ram_block1a23.port_a_byte_size = 1;
defparam ram_block1a23.port_a_data_out_clear = "none";
defparam ram_block1a23.port_a_data_out_clock = "none";
defparam ram_block1a23.port_a_data_width = 1;
defparam ram_block1a23.port_a_first_address = 0;
defparam ram_block1a23.port_a_first_bit_number = 23;
defparam ram_block1a23.port_a_last_address = 5119;
defparam ram_block1a23.port_a_logical_ram_depth = 5120;
defparam ram_block1a23.port_a_logical_ram_width = 32;
defparam ram_block1a23.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a23.ram_block_type = "auto";
defparam ram_block1a23.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a23.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a23.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a24(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[24]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a24_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a24.clk0_core_clock_enable = "ena0";
defparam ram_block1a24.clk0_input_clock_enable = "ena0";
defparam ram_block1a24.data_interleave_offset_in_bits = 1;
defparam ram_block1a24.data_interleave_width_in_bits = 1;
defparam ram_block1a24.init_file = "first_nios2_system_onchip_mem.hex";
defparam ram_block1a24.init_file_layout = "port_a";
defparam ram_block1a24.logical_ram_name = "first_nios2_system_onchip_mem:onchip_mem|altsyncram:the_altsyncram|altsyncram_mun1:auto_generated|ALTSYNCRAM";
defparam ram_block1a24.operation_mode = "single_port";
defparam ram_block1a24.port_a_address_clear = "none";
defparam ram_block1a24.port_a_address_width = 13;
defparam ram_block1a24.port_a_byte_enable_mask_width = 1;
defparam ram_block1a24.port_a_byte_size = 1;
defparam ram_block1a24.port_a_data_out_clear = "none";
defparam ram_block1a24.port_a_data_out_clock = "none";
defparam ram_block1a24.port_a_data_width = 1;
defparam ram_block1a24.port_a_first_address = 0;
defparam ram_block1a24.port_a_first_bit_number = 24;
defparam ram_block1a24.port_a_last_address = 5119;
defparam ram_block1a24.port_a_logical_ram_depth = 5120;
defparam ram_block1a24.port_a_logical_ram_width = 32;
defparam ram_block1a24.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a24.ram_block_type = "auto";
defparam ram_block1a24.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a24.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a24.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a25(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[25]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a25_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a25.clk0_core_clock_enable = "ena0";
defparam ram_block1a25.clk0_input_clock_enable = "ena0";
defparam ram_block1a25.data_interleave_offset_in_bits = 1;
defparam ram_block1a25.data_interleave_width_in_bits = 1;
defparam ram_block1a25.init_file = "first_nios2_system_onchip_mem.hex";
defparam ram_block1a25.init_file_layout = "port_a";
defparam ram_block1a25.logical_ram_name = "first_nios2_system_onchip_mem:onchip_mem|altsyncram:the_altsyncram|altsyncram_mun1:auto_generated|ALTSYNCRAM";
defparam ram_block1a25.operation_mode = "single_port";
defparam ram_block1a25.port_a_address_clear = "none";
defparam ram_block1a25.port_a_address_width = 13;
defparam ram_block1a25.port_a_byte_enable_mask_width = 1;
defparam ram_block1a25.port_a_byte_size = 1;
defparam ram_block1a25.port_a_data_out_clear = "none";
defparam ram_block1a25.port_a_data_out_clock = "none";
defparam ram_block1a25.port_a_data_width = 1;
defparam ram_block1a25.port_a_first_address = 0;
defparam ram_block1a25.port_a_first_bit_number = 25;
defparam ram_block1a25.port_a_last_address = 5119;
defparam ram_block1a25.port_a_logical_ram_depth = 5120;
defparam ram_block1a25.port_a_logical_ram_width = 32;
defparam ram_block1a25.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a25.ram_block_type = "auto";
defparam ram_block1a25.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a25.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a25.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a31(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a31_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a31.clk0_core_clock_enable = "ena0";
defparam ram_block1a31.clk0_input_clock_enable = "ena0";
defparam ram_block1a31.data_interleave_offset_in_bits = 1;
defparam ram_block1a31.data_interleave_width_in_bits = 1;
defparam ram_block1a31.init_file = "first_nios2_system_onchip_mem.hex";
defparam ram_block1a31.init_file_layout = "port_a";
defparam ram_block1a31.logical_ram_name = "first_nios2_system_onchip_mem:onchip_mem|altsyncram:the_altsyncram|altsyncram_mun1:auto_generated|ALTSYNCRAM";
defparam ram_block1a31.operation_mode = "single_port";
defparam ram_block1a31.port_a_address_clear = "none";
defparam ram_block1a31.port_a_address_width = 13;
defparam ram_block1a31.port_a_byte_enable_mask_width = 1;
defparam ram_block1a31.port_a_byte_size = 1;
defparam ram_block1a31.port_a_data_out_clear = "none";
defparam ram_block1a31.port_a_data_out_clock = "none";
defparam ram_block1a31.port_a_data_width = 1;
defparam ram_block1a31.port_a_first_address = 0;
defparam ram_block1a31.port_a_first_bit_number = 31;
defparam ram_block1a31.port_a_last_address = 5119;
defparam ram_block1a31.port_a_logical_ram_depth = 5120;
defparam ram_block1a31.port_a_logical_ram_width = 32;
defparam ram_block1a31.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a31.ram_block_type = "auto";
defparam ram_block1a31.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a31.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a31.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a21(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a21_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a21.clk0_core_clock_enable = "ena0";
defparam ram_block1a21.clk0_input_clock_enable = "ena0";
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.init_file = "first_nios2_system_onchip_mem.hex";
defparam ram_block1a21.init_file_layout = "port_a";
defparam ram_block1a21.logical_ram_name = "first_nios2_system_onchip_mem:onchip_mem|altsyncram:the_altsyncram|altsyncram_mun1:auto_generated|ALTSYNCRAM";
defparam ram_block1a21.operation_mode = "single_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 13;
defparam ram_block1a21.port_a_byte_enable_mask_width = 1;
defparam ram_block1a21.port_a_byte_size = 1;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 5119;
defparam ram_block1a21.port_a_logical_ram_depth = 5120;
defparam ram_block1a21.port_a_logical_ram_width = 32;
defparam ram_block1a21.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a21.ram_block_type = "auto";
defparam ram_block1a21.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a21.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a21.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a11(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a11_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.clk0_input_clock_enable = "ena0";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.init_file = "first_nios2_system_onchip_mem.hex";
defparam ram_block1a11.init_file_layout = "port_a";
defparam ram_block1a11.logical_ram_name = "first_nios2_system_onchip_mem:onchip_mem|altsyncram:the_altsyncram|altsyncram_mun1:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.operation_mode = "single_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 13;
defparam ram_block1a11.port_a_byte_enable_mask_width = 1;
defparam ram_block1a11.port_a_byte_size = 1;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 5119;
defparam ram_block1a11.port_a_logical_ram_depth = 5120;
defparam ram_block1a11.port_a_logical_ram_width = 32;
defparam ram_block1a11.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a11.ram_block_type = "auto";
defparam ram_block1a11.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a11.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a11.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a28(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[28]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a28_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a28.clk0_core_clock_enable = "ena0";
defparam ram_block1a28.clk0_input_clock_enable = "ena0";
defparam ram_block1a28.data_interleave_offset_in_bits = 1;
defparam ram_block1a28.data_interleave_width_in_bits = 1;
defparam ram_block1a28.init_file = "first_nios2_system_onchip_mem.hex";
defparam ram_block1a28.init_file_layout = "port_a";
defparam ram_block1a28.logical_ram_name = "first_nios2_system_onchip_mem:onchip_mem|altsyncram:the_altsyncram|altsyncram_mun1:auto_generated|ALTSYNCRAM";
defparam ram_block1a28.operation_mode = "single_port";
defparam ram_block1a28.port_a_address_clear = "none";
defparam ram_block1a28.port_a_address_width = 13;
defparam ram_block1a28.port_a_byte_enable_mask_width = 1;
defparam ram_block1a28.port_a_byte_size = 1;
defparam ram_block1a28.port_a_data_out_clear = "none";
defparam ram_block1a28.port_a_data_out_clock = "none";
defparam ram_block1a28.port_a_data_width = 1;
defparam ram_block1a28.port_a_first_address = 0;
defparam ram_block1a28.port_a_first_bit_number = 28;
defparam ram_block1a28.port_a_last_address = 5119;
defparam ram_block1a28.port_a_logical_ram_depth = 5120;
defparam ram_block1a28.port_a_logical_ram_width = 32;
defparam ram_block1a28.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a28.ram_block_type = "auto";
defparam ram_block1a28.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a28.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a28.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a10(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a10_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.clk0_input_clock_enable = "ena0";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.init_file = "first_nios2_system_onchip_mem.hex";
defparam ram_block1a10.init_file_layout = "port_a";
defparam ram_block1a10.logical_ram_name = "first_nios2_system_onchip_mem:onchip_mem|altsyncram:the_altsyncram|altsyncram_mun1:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.operation_mode = "single_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 13;
defparam ram_block1a10.port_a_byte_enable_mask_width = 1;
defparam ram_block1a10.port_a_byte_size = 1;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 5119;
defparam ram_block1a10.port_a_logical_ram_depth = 5120;
defparam ram_block1a10.port_a_logical_ram_width = 32;
defparam ram_block1a10.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a10.ram_block_type = "auto";
defparam ram_block1a10.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a10.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a10.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a27(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[27]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a27_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a27.clk0_core_clock_enable = "ena0";
defparam ram_block1a27.clk0_input_clock_enable = "ena0";
defparam ram_block1a27.data_interleave_offset_in_bits = 1;
defparam ram_block1a27.data_interleave_width_in_bits = 1;
defparam ram_block1a27.init_file = "first_nios2_system_onchip_mem.hex";
defparam ram_block1a27.init_file_layout = "port_a";
defparam ram_block1a27.logical_ram_name = "first_nios2_system_onchip_mem:onchip_mem|altsyncram:the_altsyncram|altsyncram_mun1:auto_generated|ALTSYNCRAM";
defparam ram_block1a27.operation_mode = "single_port";
defparam ram_block1a27.port_a_address_clear = "none";
defparam ram_block1a27.port_a_address_width = 13;
defparam ram_block1a27.port_a_byte_enable_mask_width = 1;
defparam ram_block1a27.port_a_byte_size = 1;
defparam ram_block1a27.port_a_data_out_clear = "none";
defparam ram_block1a27.port_a_data_out_clock = "none";
defparam ram_block1a27.port_a_data_width = 1;
defparam ram_block1a27.port_a_first_address = 0;
defparam ram_block1a27.port_a_first_bit_number = 27;
defparam ram_block1a27.port_a_last_address = 5119;
defparam ram_block1a27.port_a_logical_ram_depth = 5120;
defparam ram_block1a27.port_a_logical_ram_width = 32;
defparam ram_block1a27.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a27.ram_block_type = "auto";
defparam ram_block1a27.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a27.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a27.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a8(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a8_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk0_input_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.init_file = "first_nios2_system_onchip_mem.hex";
defparam ram_block1a8.init_file_layout = "port_a";
defparam ram_block1a8.logical_ram_name = "first_nios2_system_onchip_mem:onchip_mem|altsyncram:the_altsyncram|altsyncram_mun1:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.operation_mode = "single_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 13;
defparam ram_block1a8.port_a_byte_enable_mask_width = 1;
defparam ram_block1a8.port_a_byte_size = 1;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 5119;
defparam ram_block1a8.port_a_logical_ram_depth = 5120;
defparam ram_block1a8.port_a_logical_ram_width = 32;
defparam ram_block1a8.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a8.ram_block_type = "auto";
defparam ram_block1a8.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a8.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a8.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a9(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a9_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk0_input_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.init_file = "first_nios2_system_onchip_mem.hex";
defparam ram_block1a9.init_file_layout = "port_a";
defparam ram_block1a9.logical_ram_name = "first_nios2_system_onchip_mem:onchip_mem|altsyncram:the_altsyncram|altsyncram_mun1:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.operation_mode = "single_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 13;
defparam ram_block1a9.port_a_byte_enable_mask_width = 1;
defparam ram_block1a9.port_a_byte_size = 1;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 5119;
defparam ram_block1a9.port_a_logical_ram_depth = 5120;
defparam ram_block1a9.port_a_logical_ram_width = 32;
defparam ram_block1a9.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a9.ram_block_type = "auto";
defparam ram_block1a9.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a9.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a9.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a26(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[26]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a26_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a26.clk0_core_clock_enable = "ena0";
defparam ram_block1a26.clk0_input_clock_enable = "ena0";
defparam ram_block1a26.data_interleave_offset_in_bits = 1;
defparam ram_block1a26.data_interleave_width_in_bits = 1;
defparam ram_block1a26.init_file = "first_nios2_system_onchip_mem.hex";
defparam ram_block1a26.init_file_layout = "port_a";
defparam ram_block1a26.logical_ram_name = "first_nios2_system_onchip_mem:onchip_mem|altsyncram:the_altsyncram|altsyncram_mun1:auto_generated|ALTSYNCRAM";
defparam ram_block1a26.operation_mode = "single_port";
defparam ram_block1a26.port_a_address_clear = "none";
defparam ram_block1a26.port_a_address_width = 13;
defparam ram_block1a26.port_a_byte_enable_mask_width = 1;
defparam ram_block1a26.port_a_byte_size = 1;
defparam ram_block1a26.port_a_data_out_clear = "none";
defparam ram_block1a26.port_a_data_out_clock = "none";
defparam ram_block1a26.port_a_data_width = 1;
defparam ram_block1a26.port_a_first_address = 0;
defparam ram_block1a26.port_a_first_bit_number = 26;
defparam ram_block1a26.port_a_last_address = 5119;
defparam ram_block1a26.port_a_logical_ram_depth = 5120;
defparam ram_block1a26.port_a_logical_ram_width = 32;
defparam ram_block1a26.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a26.ram_block_type = "auto";
defparam ram_block1a26.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a26.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a26.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a20(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a20_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a20.clk0_core_clock_enable = "ena0";
defparam ram_block1a20.clk0_input_clock_enable = "ena0";
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.init_file = "first_nios2_system_onchip_mem.hex";
defparam ram_block1a20.init_file_layout = "port_a";
defparam ram_block1a20.logical_ram_name = "first_nios2_system_onchip_mem:onchip_mem|altsyncram:the_altsyncram|altsyncram_mun1:auto_generated|ALTSYNCRAM";
defparam ram_block1a20.operation_mode = "single_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 13;
defparam ram_block1a20.port_a_byte_enable_mask_width = 1;
defparam ram_block1a20.port_a_byte_size = 1;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 5119;
defparam ram_block1a20.port_a_logical_ram_depth = 5120;
defparam ram_block1a20.port_a_logical_ram_width = 32;
defparam ram_block1a20.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a20.ram_block_type = "auto";
defparam ram_block1a20.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a20.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a20.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a19(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a19_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a19.clk0_core_clock_enable = "ena0";
defparam ram_block1a19.clk0_input_clock_enable = "ena0";
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.init_file = "first_nios2_system_onchip_mem.hex";
defparam ram_block1a19.init_file_layout = "port_a";
defparam ram_block1a19.logical_ram_name = "first_nios2_system_onchip_mem:onchip_mem|altsyncram:the_altsyncram|altsyncram_mun1:auto_generated|ALTSYNCRAM";
defparam ram_block1a19.operation_mode = "single_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 13;
defparam ram_block1a19.port_a_byte_enable_mask_width = 1;
defparam ram_block1a19.port_a_byte_size = 1;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 5119;
defparam ram_block1a19.port_a_logical_ram_depth = 5120;
defparam ram_block1a19.port_a_logical_ram_width = 32;
defparam ram_block1a19.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a19.ram_block_type = "auto";
defparam ram_block1a19.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a19.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a19.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a17(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a17_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a17.clk0_core_clock_enable = "ena0";
defparam ram_block1a17.clk0_input_clock_enable = "ena0";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.init_file = "first_nios2_system_onchip_mem.hex";
defparam ram_block1a17.init_file_layout = "port_a";
defparam ram_block1a17.logical_ram_name = "first_nios2_system_onchip_mem:onchip_mem|altsyncram:the_altsyncram|altsyncram_mun1:auto_generated|ALTSYNCRAM";
defparam ram_block1a17.operation_mode = "single_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 13;
defparam ram_block1a17.port_a_byte_enable_mask_width = 1;
defparam ram_block1a17.port_a_byte_size = 1;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 5119;
defparam ram_block1a17.port_a_logical_ram_depth = 5120;
defparam ram_block1a17.port_a_logical_ram_width = 32;
defparam ram_block1a17.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a17.ram_block_type = "auto";
defparam ram_block1a17.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a17.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a17.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a30(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[30]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a30_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a30.clk0_core_clock_enable = "ena0";
defparam ram_block1a30.clk0_input_clock_enable = "ena0";
defparam ram_block1a30.data_interleave_offset_in_bits = 1;
defparam ram_block1a30.data_interleave_width_in_bits = 1;
defparam ram_block1a30.init_file = "first_nios2_system_onchip_mem.hex";
defparam ram_block1a30.init_file_layout = "port_a";
defparam ram_block1a30.logical_ram_name = "first_nios2_system_onchip_mem:onchip_mem|altsyncram:the_altsyncram|altsyncram_mun1:auto_generated|ALTSYNCRAM";
defparam ram_block1a30.operation_mode = "single_port";
defparam ram_block1a30.port_a_address_clear = "none";
defparam ram_block1a30.port_a_address_width = 13;
defparam ram_block1a30.port_a_byte_enable_mask_width = 1;
defparam ram_block1a30.port_a_byte_size = 1;
defparam ram_block1a30.port_a_data_out_clear = "none";
defparam ram_block1a30.port_a_data_out_clock = "none";
defparam ram_block1a30.port_a_data_width = 1;
defparam ram_block1a30.port_a_first_address = 0;
defparam ram_block1a30.port_a_first_bit_number = 30;
defparam ram_block1a30.port_a_last_address = 5119;
defparam ram_block1a30.port_a_logical_ram_depth = 5120;
defparam ram_block1a30.port_a_logical_ram_width = 32;
defparam ram_block1a30.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a30.ram_block_type = "auto";
defparam ram_block1a30.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a30.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a30.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a18(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a18_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a18.clk0_core_clock_enable = "ena0";
defparam ram_block1a18.clk0_input_clock_enable = "ena0";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.init_file = "first_nios2_system_onchip_mem.hex";
defparam ram_block1a18.init_file_layout = "port_a";
defparam ram_block1a18.logical_ram_name = "first_nios2_system_onchip_mem:onchip_mem|altsyncram:the_altsyncram|altsyncram_mun1:auto_generated|ALTSYNCRAM";
defparam ram_block1a18.operation_mode = "single_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 13;
defparam ram_block1a18.port_a_byte_enable_mask_width = 1;
defparam ram_block1a18.port_a_byte_size = 1;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 5119;
defparam ram_block1a18.port_a_logical_ram_depth = 5120;
defparam ram_block1a18.port_a_logical_ram_width = 32;
defparam ram_block1a18.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a18.ram_block_type = "auto";
defparam ram_block1a18.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a18.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a18.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a16(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a16_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a16.clk0_core_clock_enable = "ena0";
defparam ram_block1a16.clk0_input_clock_enable = "ena0";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.init_file = "first_nios2_system_onchip_mem.hex";
defparam ram_block1a16.init_file_layout = "port_a";
defparam ram_block1a16.logical_ram_name = "first_nios2_system_onchip_mem:onchip_mem|altsyncram:the_altsyncram|altsyncram_mun1:auto_generated|ALTSYNCRAM";
defparam ram_block1a16.operation_mode = "single_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 13;
defparam ram_block1a16.port_a_byte_enable_mask_width = 1;
defparam ram_block1a16.port_a_byte_size = 1;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 5119;
defparam ram_block1a16.port_a_logical_ram_depth = 5120;
defparam ram_block1a16.port_a_logical_ram_width = 32;
defparam ram_block1a16.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a16.ram_block_type = "auto";
defparam ram_block1a16.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a16.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a16.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a15(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a15_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.clk0_input_clock_enable = "ena0";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.init_file = "first_nios2_system_onchip_mem.hex";
defparam ram_block1a15.init_file_layout = "port_a";
defparam ram_block1a15.logical_ram_name = "first_nios2_system_onchip_mem:onchip_mem|altsyncram:the_altsyncram|altsyncram_mun1:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.operation_mode = "single_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 13;
defparam ram_block1a15.port_a_byte_enable_mask_width = 1;
defparam ram_block1a15.port_a_byte_size = 1;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 5119;
defparam ram_block1a15.port_a_logical_ram_depth = 5120;
defparam ram_block1a15.port_a_logical_ram_width = 32;
defparam ram_block1a15.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a15.ram_block_type = "auto";
defparam ram_block1a15.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a15.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a15.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a12(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a12_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.clk0_input_clock_enable = "ena0";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.init_file = "first_nios2_system_onchip_mem.hex";
defparam ram_block1a12.init_file_layout = "port_a";
defparam ram_block1a12.logical_ram_name = "first_nios2_system_onchip_mem:onchip_mem|altsyncram:the_altsyncram|altsyncram_mun1:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.operation_mode = "single_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 13;
defparam ram_block1a12.port_a_byte_enable_mask_width = 1;
defparam ram_block1a12.port_a_byte_size = 1;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 5119;
defparam ram_block1a12.port_a_logical_ram_depth = 5120;
defparam ram_block1a12.port_a_logical_ram_width = 32;
defparam ram_block1a12.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a12.ram_block_type = "auto";
defparam ram_block1a12.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a12.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a12.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a13(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a13_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.clk0_input_clock_enable = "ena0";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.init_file = "first_nios2_system_onchip_mem.hex";
defparam ram_block1a13.init_file_layout = "port_a";
defparam ram_block1a13.logical_ram_name = "first_nios2_system_onchip_mem:onchip_mem|altsyncram:the_altsyncram|altsyncram_mun1:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.operation_mode = "single_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 13;
defparam ram_block1a13.port_a_byte_enable_mask_width = 1;
defparam ram_block1a13.port_a_byte_size = 1;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 5119;
defparam ram_block1a13.port_a_logical_ram_depth = 5120;
defparam ram_block1a13.port_a_logical_ram_width = 32;
defparam ram_block1a13.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a13.ram_block_type = "auto";
defparam ram_block1a13.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a13.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a13.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a14(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a14_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.clk0_input_clock_enable = "ena0";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.init_file = "first_nios2_system_onchip_mem.hex";
defparam ram_block1a14.init_file_layout = "port_a";
defparam ram_block1a14.logical_ram_name = "first_nios2_system_onchip_mem:onchip_mem|altsyncram:the_altsyncram|altsyncram_mun1:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.operation_mode = "single_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 13;
defparam ram_block1a14.port_a_byte_enable_mask_width = 1;
defparam ram_block1a14.port_a_byte_size = 1;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 5119;
defparam ram_block1a14.port_a_logical_ram_depth = 5120;
defparam ram_block1a14.port_a_logical_ram_width = 32;
defparam ram_block1a14.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a14.ram_block_type = "auto";
defparam ram_block1a14.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a14.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a14.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a29(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[29]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a29_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a29.clk0_core_clock_enable = "ena0";
defparam ram_block1a29.clk0_input_clock_enable = "ena0";
defparam ram_block1a29.data_interleave_offset_in_bits = 1;
defparam ram_block1a29.data_interleave_width_in_bits = 1;
defparam ram_block1a29.init_file = "first_nios2_system_onchip_mem.hex";
defparam ram_block1a29.init_file_layout = "port_a";
defparam ram_block1a29.logical_ram_name = "first_nios2_system_onchip_mem:onchip_mem|altsyncram:the_altsyncram|altsyncram_mun1:auto_generated|ALTSYNCRAM";
defparam ram_block1a29.operation_mode = "single_port";
defparam ram_block1a29.port_a_address_clear = "none";
defparam ram_block1a29.port_a_address_width = 13;
defparam ram_block1a29.port_a_byte_enable_mask_width = 1;
defparam ram_block1a29.port_a_byte_size = 1;
defparam ram_block1a29.port_a_data_out_clear = "none";
defparam ram_block1a29.port_a_data_out_clock = "none";
defparam ram_block1a29.port_a_data_width = 1;
defparam ram_block1a29.port_a_first_address = 0;
defparam ram_block1a29.port_a_first_bit_number = 29;
defparam ram_block1a29.port_a_last_address = 5119;
defparam ram_block1a29.port_a_logical_ram_depth = 5120;
defparam ram_block1a29.port_a_logical_ram_width = 32;
defparam ram_block1a29.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a29.ram_block_type = "auto";
defparam ram_block1a29.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a29.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a29.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

endmodule

module first_nios2_system_first_nios2_system_rtd1 (
	readdata_0,
	Equal0,
	r_sync_rst,
	clk_clk,
	rtd1_external_connection_export)/* synthesis synthesis_greybox=1 */;
output 	readdata_0;
input 	Equal0;
input 	r_sync_rst;
input 	clk_clk;
input 	rtd1_external_connection_export;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \readdata[0] (
	.clk(clk_clk),
	.d(rtd1_external_connection_export),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(Equal0),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_0),
	.prn(vcc));
defparam \readdata[0] .is_wysiwyg = "true";
defparam \readdata[0] .power_up = "low";

endmodule

module first_nios2_system_first_nios2_system_rtd1_1 (
	readdata_0,
	Equal0,
	r_sync_rst,
	clk_clk,
	rtd2_external_connection_export)/* synthesis synthesis_greybox=1 */;
output 	readdata_0;
input 	Equal0;
input 	r_sync_rst;
input 	clk_clk;
input 	rtd2_external_connection_export;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \readdata[0] (
	.clk(clk_clk),
	.d(rtd2_external_connection_export),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(Equal0),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_0),
	.prn(vcc));
defparam \readdata[0] .is_wysiwyg = "true";
defparam \readdata[0] .power_up = "low";

endmodule

module first_nios2_system_first_nios2_system_sys_clk_timer (
	writedata,
	A_mem_baddr_4,
	clr_break_line,
	d_write,
	A_mem_baddr_3,
	A_mem_baddr_2,
	reset_n,
	Equal2,
	wait_latency_counter_0,
	mem_used_1,
	wait_latency_counter_1,
	timeout_occurred1,
	control_register_0,
	readdata_0,
	readdata_1,
	readdata_2,
	readdata_3,
	readdata_4,
	readdata_5,
	readdata_6,
	readdata_7,
	readdata_11,
	readdata_10,
	readdata_8,
	readdata_9,
	readdata_15,
	readdata_12,
	readdata_13,
	readdata_14,
	clk)/* synthesis synthesis_greybox=1 */;
input 	[15:0] writedata;
input 	A_mem_baddr_4;
input 	clr_break_line;
input 	d_write;
input 	A_mem_baddr_3;
input 	A_mem_baddr_2;
input 	reset_n;
input 	Equal2;
input 	wait_latency_counter_0;
input 	mem_used_1;
input 	wait_latency_counter_1;
output 	timeout_occurred1;
output 	control_register_0;
output 	readdata_0;
output 	readdata_1;
output 	readdata_2;
output 	readdata_3;
output 	readdata_4;
output 	readdata_5;
output 	readdata_6;
output 	readdata_7;
output 	readdata_11;
output 	readdata_10;
output 	readdata_8;
output 	readdata_9;
output 	readdata_15;
output 	readdata_12;
output 	readdata_13;
output 	readdata_14;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \period_l_wr_strobe~0_combout ;
wire \period_l_wr_strobe~1_combout ;
wire \status_wr_strobe~0_combout ;
wire \period_l_register[6]~5_combout ;
wire \Equal6~2_combout ;
wire \period_l_wr_strobe~combout ;
wire \period_l_register[6]~q ;
wire \period_l_register[3]~0_combout ;
wire \period_l_register[3]~q ;
wire \period_l_register[2]~6_combout ;
wire \period_l_register[2]~q ;
wire \period_l_register[1]~7_combout ;
wire \period_l_register[1]~q ;
wire \period_l_register[0]~8_combout ;
wire \period_l_register[0]~q ;
wire \Add0~117_sumout ;
wire \internal_counter~8_combout ;
wire \force_reload~0_combout ;
wire \force_reload~q ;
wire \Equal6~0_combout ;
wire \control_wr_strobe~combout ;
wire \control_register[1]~q ;
wire \counter_is_running~0_combout ;
wire \counter_is_running~1_combout ;
wire \counter_is_running~q ;
wire \always0~1_combout ;
wire \internal_counter[0]~q ;
wire \Add0~118 ;
wire \Add0~113_sumout ;
wire \internal_counter~7_combout ;
wire \internal_counter[1]~q ;
wire \Add0~114 ;
wire \Add0~109_sumout ;
wire \internal_counter~6_combout ;
wire \internal_counter[2]~q ;
wire \Add0~110 ;
wire \Add0~57_sumout ;
wire \internal_counter~0_combout ;
wire \internal_counter[3]~q ;
wire \Add0~58 ;
wire \Add0~125_sumout ;
wire \period_l_register[4]~q ;
wire \internal_counter[4]~q ;
wire \Add0~126 ;
wire \Add0~121_sumout ;
wire \period_l_register[5]~q ;
wire \internal_counter[5]~q ;
wire \Add0~122 ;
wire \Add0~105_sumout ;
wire \internal_counter~5_combout ;
wire \internal_counter[6]~q ;
wire \Add0~106 ;
wire \Add0~5_sumout ;
wire \period_l_register[7]~q ;
wire \internal_counter[7]~q ;
wire \period_l_register[15]~1_combout ;
wire \period_l_register[15]~q ;
wire \period_l_register[14]~2_combout ;
wire \period_l_register[14]~q ;
wire \Add0~2 ;
wire \Add0~29_sumout ;
wire \period_l_register[11]~q ;
wire \internal_counter[11]~q ;
wire \Add0~30 ;
wire \Add0~25_sumout ;
wire \period_l_register[12]~q ;
wire \internal_counter[12]~q ;
wire \Add0~26 ;
wire \Add0~21_sumout ;
wire \period_l_register[13]~q ;
wire \internal_counter[13]~q ;
wire \Add0~22 ;
wire \Add0~93_sumout ;
wire \internal_counter~2_combout ;
wire \internal_counter[14]~q ;
wire \Add0~94 ;
wire \Add0~89_sumout ;
wire \internal_counter~1_combout ;
wire \internal_counter[15]~q ;
wire \Add0~90 ;
wire \Add0~17_sumout ;
wire \Equal6~1_combout ;
wire \period_h_wr_strobe~combout ;
wire \period_h_register[0]~q ;
wire \internal_counter[16]~q ;
wire \Add0~18 ;
wire \Add0~13_sumout ;
wire \period_h_register[1]~q ;
wire \internal_counter[17]~q ;
wire \Add0~14 ;
wire \Add0~9_sumout ;
wire \period_h_register[2]~q ;
wire \internal_counter[18]~q ;
wire \Equal0~0_combout ;
wire \Add0~10 ;
wire \Add0~53_sumout ;
wire \period_h_register[3]~q ;
wire \internal_counter[19]~q ;
wire \Add0~54 ;
wire \Add0~61_sumout ;
wire \period_h_register[4]~q ;
wire \internal_counter[20]~q ;
wire \Add0~62 ;
wire \Add0~49_sumout ;
wire \period_h_register[5]~q ;
wire \internal_counter[21]~q ;
wire \Add0~50 ;
wire \Add0~45_sumout ;
wire \period_h_register[6]~q ;
wire \internal_counter[22]~q ;
wire \Add0~46 ;
wire \Add0~41_sumout ;
wire \period_h_register[7]~q ;
wire \internal_counter[23]~q ;
wire \Add0~42 ;
wire \Add0~69_sumout ;
wire \period_h_register[8]~q ;
wire \internal_counter[24]~q ;
wire \Add0~70 ;
wire \Add0~37_sumout ;
wire \period_h_register[9]~q ;
wire \internal_counter[25]~q ;
wire \Add0~38 ;
wire \Add0~33_sumout ;
wire \period_h_register[10]~q ;
wire \internal_counter[26]~q ;
wire \Equal0~1_combout ;
wire \Add0~34 ;
wire \Add0~65_sumout ;
wire \period_h_register[11]~q ;
wire \internal_counter[27]~q ;
wire \Add0~66 ;
wire \Add0~85_sumout ;
wire \period_h_register[12]~q ;
wire \internal_counter[28]~q ;
wire \Add0~86 ;
wire \Add0~81_sumout ;
wire \period_h_register[13]~q ;
wire \internal_counter[29]~q ;
wire \Add0~82 ;
wire \Add0~77_sumout ;
wire \period_h_register[14]~q ;
wire \internal_counter[30]~q ;
wire \Add0~78 ;
wire \Add0~73_sumout ;
wire \period_h_register[15]~q ;
wire \internal_counter[31]~q ;
wire \Equal0~2_combout ;
wire \period_l_register[8]~4_combout ;
wire \period_l_register[8]~q ;
wire \Add0~6 ;
wire \Add0~101_sumout ;
wire \internal_counter~4_combout ;
wire \internal_counter[8]~q ;
wire \Equal0~3_combout ;
wire \Equal0~4_combout ;
wire \Equal0~5_combout ;
wire \always0~0_combout ;
wire \period_l_register[9]~3_combout ;
wire \period_l_register[9]~q ;
wire \Add0~102 ;
wire \Add0~97_sumout ;
wire \internal_counter~3_combout ;
wire \internal_counter[9]~q ;
wire \Add0~98 ;
wire \Add0~1_sumout ;
wire \period_l_register[10]~q ;
wire \internal_counter[10]~q ;
wire \Equal0~6_combout ;
wire \delayed_unxcounter_is_zeroxx0~q ;
wire \timeout_occurred~0_combout ;
wire \counter_snapshot[0]~0_combout ;
wire \Equal6~3_combout ;
wire \snap_strobe~0_combout ;
wire \counter_snapshot[0]~q ;
wire \Equal6~4_combout ;
wire \read_mux_out[0]~0_combout ;
wire \counter_snapshot[16]~q ;
wire \read_mux_out[0]~1_combout ;
wire \read_mux_out[0]~combout ;
wire \counter_snapshot[1]~1_combout ;
wire \counter_snapshot[1]~q ;
wire \read_mux_out[1]~2_combout ;
wire \counter_snapshot[17]~q ;
wire \read_mux_out[1]~3_combout ;
wire \read_mux_out[1]~combout ;
wire \counter_snapshot[2]~2_combout ;
wire \counter_snapshot[2]~q ;
wire \read_mux_out[2]~4_combout ;
wire \Equal6~5_combout ;
wire \counter_snapshot[18]~q ;
wire \control_register[2]~q ;
wire \read_mux_out[2]~5_combout ;
wire \read_mux_out[2]~combout ;
wire \counter_snapshot[3]~3_combout ;
wire \counter_snapshot[3]~q ;
wire \read_mux_out[3]~6_combout ;
wire \counter_snapshot[19]~q ;
wire \control_register[3]~q ;
wire \read_mux_out[3]~7_combout ;
wire \read_mux_out[3]~combout ;
wire \counter_snapshot[4]~q ;
wire \counter_snapshot[20]~q ;
wire \read_mux_out[4]~52_combout ;
wire \counter_snapshot[5]~q ;
wire \counter_snapshot[21]~q ;
wire \read_mux_out[5]~48_combout ;
wire \counter_snapshot[6]~4_combout ;
wire \counter_snapshot[6]~q ;
wire \counter_snapshot[22]~q ;
wire \read_mux_out[6]~44_combout ;
wire \counter_snapshot[7]~q ;
wire \counter_snapshot[23]~q ;
wire \read_mux_out[7]~40_combout ;
wire \counter_snapshot[11]~q ;
wire \counter_snapshot[27]~q ;
wire \read_mux_out[11]~36_combout ;
wire \counter_snapshot[10]~q ;
wire \counter_snapshot[26]~q ;
wire \read_mux_out[10]~32_combout ;
wire \counter_snapshot[8]~5_combout ;
wire \counter_snapshot[8]~q ;
wire \counter_snapshot[24]~q ;
wire \read_mux_out[8]~28_combout ;
wire \counter_snapshot[9]~6_combout ;
wire \counter_snapshot[9]~q ;
wire \counter_snapshot[25]~q ;
wire \read_mux_out[9]~24_combout ;
wire \counter_snapshot[15]~7_combout ;
wire \counter_snapshot[15]~q ;
wire \counter_snapshot[31]~q ;
wire \read_mux_out[15]~20_combout ;
wire \counter_snapshot[12]~q ;
wire \counter_snapshot[28]~q ;
wire \read_mux_out[12]~16_combout ;
wire \counter_snapshot[13]~q ;
wire \counter_snapshot[29]~q ;
wire \read_mux_out[13]~12_combout ;
wire \counter_snapshot[14]~8_combout ;
wire \counter_snapshot[14]~q ;
wire \counter_snapshot[30]~q ;
wire \read_mux_out[14]~8_combout ;


dffeas timeout_occurred(
	.clk(clk),
	.d(\timeout_occurred~0_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(timeout_occurred1),
	.prn(vcc));
defparam timeout_occurred.is_wysiwyg = "true";
defparam timeout_occurred.power_up = "low";

dffeas \control_register[0] (
	.clk(clk),
	.d(writedata[0]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\control_wr_strobe~combout ),
	.q(control_register_0),
	.prn(vcc));
defparam \control_register[0] .is_wysiwyg = "true";
defparam \control_register[0] .power_up = "low";

dffeas \readdata[0] (
	.clk(clk),
	.d(\read_mux_out[0]~combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_0),
	.prn(vcc));
defparam \readdata[0] .is_wysiwyg = "true";
defparam \readdata[0] .power_up = "low";

dffeas \readdata[1] (
	.clk(clk),
	.d(\read_mux_out[1]~combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_1),
	.prn(vcc));
defparam \readdata[1] .is_wysiwyg = "true";
defparam \readdata[1] .power_up = "low";

dffeas \readdata[2] (
	.clk(clk),
	.d(\read_mux_out[2]~combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_2),
	.prn(vcc));
defparam \readdata[2] .is_wysiwyg = "true";
defparam \readdata[2] .power_up = "low";

dffeas \readdata[3] (
	.clk(clk),
	.d(\read_mux_out[3]~combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_3),
	.prn(vcc));
defparam \readdata[3] .is_wysiwyg = "true";
defparam \readdata[3] .power_up = "low";

dffeas \readdata[4] (
	.clk(clk),
	.d(\read_mux_out[4]~52_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_4),
	.prn(vcc));
defparam \readdata[4] .is_wysiwyg = "true";
defparam \readdata[4] .power_up = "low";

dffeas \readdata[5] (
	.clk(clk),
	.d(\read_mux_out[5]~48_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_5),
	.prn(vcc));
defparam \readdata[5] .is_wysiwyg = "true";
defparam \readdata[5] .power_up = "low";

dffeas \readdata[6] (
	.clk(clk),
	.d(\read_mux_out[6]~44_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_6),
	.prn(vcc));
defparam \readdata[6] .is_wysiwyg = "true";
defparam \readdata[6] .power_up = "low";

dffeas \readdata[7] (
	.clk(clk),
	.d(\read_mux_out[7]~40_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_7),
	.prn(vcc));
defparam \readdata[7] .is_wysiwyg = "true";
defparam \readdata[7] .power_up = "low";

dffeas \readdata[11] (
	.clk(clk),
	.d(\read_mux_out[11]~36_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_11),
	.prn(vcc));
defparam \readdata[11] .is_wysiwyg = "true";
defparam \readdata[11] .power_up = "low";

dffeas \readdata[10] (
	.clk(clk),
	.d(\read_mux_out[10]~32_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_10),
	.prn(vcc));
defparam \readdata[10] .is_wysiwyg = "true";
defparam \readdata[10] .power_up = "low";

dffeas \readdata[8] (
	.clk(clk),
	.d(\read_mux_out[8]~28_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_8),
	.prn(vcc));
defparam \readdata[8] .is_wysiwyg = "true";
defparam \readdata[8] .power_up = "low";

dffeas \readdata[9] (
	.clk(clk),
	.d(\read_mux_out[9]~24_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_9),
	.prn(vcc));
defparam \readdata[9] .is_wysiwyg = "true";
defparam \readdata[9] .power_up = "low";

dffeas \readdata[15] (
	.clk(clk),
	.d(\read_mux_out[15]~20_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_15),
	.prn(vcc));
defparam \readdata[15] .is_wysiwyg = "true";
defparam \readdata[15] .power_up = "low";

dffeas \readdata[12] (
	.clk(clk),
	.d(\read_mux_out[12]~16_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_12),
	.prn(vcc));
defparam \readdata[12] .is_wysiwyg = "true";
defparam \readdata[12] .power_up = "low";

dffeas \readdata[13] (
	.clk(clk),
	.d(\read_mux_out[13]~12_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_13),
	.prn(vcc));
defparam \readdata[13] .is_wysiwyg = "true";
defparam \readdata[13] .power_up = "low";

dffeas \readdata[14] (
	.clk(clk),
	.d(\read_mux_out[14]~8_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_14),
	.prn(vcc));
defparam \readdata[14] .is_wysiwyg = "true";
defparam \readdata[14] .power_up = "low";

cyclonev_lcell_comb \period_l_wr_strobe~0 (
	.dataa(!d_write),
	.datab(!wait_latency_counter_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\period_l_wr_strobe~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \period_l_wr_strobe~0 .extended_lut = "off";
defparam \period_l_wr_strobe~0 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \period_l_wr_strobe~0 .shared_arith = "off";

cyclonev_lcell_comb \period_l_wr_strobe~1 (
	.dataa(!clr_break_line),
	.datab(!Equal2),
	.datac(!mem_used_1),
	.datad(!wait_latency_counter_1),
	.datae(!\period_l_wr_strobe~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\period_l_wr_strobe~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \period_l_wr_strobe~1 .extended_lut = "off";
defparam \period_l_wr_strobe~1 .lut_mask = 64'hFFF7FFFFFFF7FFFF;
defparam \period_l_wr_strobe~1 .shared_arith = "off";

cyclonev_lcell_comb \status_wr_strobe~0 (
	.dataa(!A_mem_baddr_3),
	.datab(!A_mem_baddr_2),
	.datac(!A_mem_baddr_4),
	.datad(!\period_l_wr_strobe~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\status_wr_strobe~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \status_wr_strobe~0 .extended_lut = "off";
defparam \status_wr_strobe~0 .lut_mask = 64'hFEFFFEFFFEFFFEFF;
defparam \status_wr_strobe~0 .shared_arith = "off";

cyclonev_lcell_comb \period_l_register[6]~5 (
	.dataa(!writedata[6]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\period_l_register[6]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \period_l_register[6]~5 .extended_lut = "off";
defparam \period_l_register[6]~5 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \period_l_register[6]~5 .shared_arith = "off";

cyclonev_lcell_comb \Equal6~2 (
	.dataa(!A_mem_baddr_3),
	.datab(!A_mem_baddr_2),
	.datac(!A_mem_baddr_4),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal6~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal6~2 .extended_lut = "off";
defparam \Equal6~2 .lut_mask = 64'hFDFDFDFDFDFDFDFD;
defparam \Equal6~2 .shared_arith = "off";

cyclonev_lcell_comb period_l_wr_strobe(
	.dataa(!clr_break_line),
	.datab(!Equal2),
	.datac(!mem_used_1),
	.datad(!wait_latency_counter_1),
	.datae(!\period_l_wr_strobe~0_combout ),
	.dataf(!\Equal6~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\period_l_wr_strobe~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam period_l_wr_strobe.extended_lut = "off";
defparam period_l_wr_strobe.lut_mask = 64'hFFF7FFFFFFFFFFFF;
defparam period_l_wr_strobe.shared_arith = "off";

dffeas \period_l_register[6] (
	.clk(clk),
	.d(\period_l_register[6]~5_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_l_wr_strobe~combout ),
	.q(\period_l_register[6]~q ),
	.prn(vcc));
defparam \period_l_register[6] .is_wysiwyg = "true";
defparam \period_l_register[6] .power_up = "low";

cyclonev_lcell_comb \period_l_register[3]~0 (
	.dataa(!writedata[3]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\period_l_register[3]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \period_l_register[3]~0 .extended_lut = "off";
defparam \period_l_register[3]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \period_l_register[3]~0 .shared_arith = "off";

dffeas \period_l_register[3] (
	.clk(clk),
	.d(\period_l_register[3]~0_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_l_wr_strobe~combout ),
	.q(\period_l_register[3]~q ),
	.prn(vcc));
defparam \period_l_register[3] .is_wysiwyg = "true";
defparam \period_l_register[3] .power_up = "low";

cyclonev_lcell_comb \period_l_register[2]~6 (
	.dataa(!writedata[2]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\period_l_register[2]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \period_l_register[2]~6 .extended_lut = "off";
defparam \period_l_register[2]~6 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \period_l_register[2]~6 .shared_arith = "off";

dffeas \period_l_register[2] (
	.clk(clk),
	.d(\period_l_register[2]~6_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_l_wr_strobe~combout ),
	.q(\period_l_register[2]~q ),
	.prn(vcc));
defparam \period_l_register[2] .is_wysiwyg = "true";
defparam \period_l_register[2] .power_up = "low";

cyclonev_lcell_comb \period_l_register[1]~7 (
	.dataa(!writedata[1]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\period_l_register[1]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \period_l_register[1]~7 .extended_lut = "off";
defparam \period_l_register[1]~7 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \period_l_register[1]~7 .shared_arith = "off";

dffeas \period_l_register[1] (
	.clk(clk),
	.d(\period_l_register[1]~7_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_l_wr_strobe~combout ),
	.q(\period_l_register[1]~q ),
	.prn(vcc));
defparam \period_l_register[1] .is_wysiwyg = "true";
defparam \period_l_register[1] .power_up = "low";

cyclonev_lcell_comb \period_l_register[0]~8 (
	.dataa(!writedata[0]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\period_l_register[0]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \period_l_register[0]~8 .extended_lut = "off";
defparam \period_l_register[0]~8 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \period_l_register[0]~8 .shared_arith = "off";

dffeas \period_l_register[0] (
	.clk(clk),
	.d(\period_l_register[0]~8_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_l_wr_strobe~combout ),
	.q(\period_l_register[0]~q ),
	.prn(vcc));
defparam \period_l_register[0] .is_wysiwyg = "true";
defparam \period_l_register[0] .power_up = "low";

cyclonev_lcell_comb \Add0~117 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\internal_counter[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~117_sumout ),
	.cout(\Add0~118 ),
	.shareout());
defparam \Add0~117 .extended_lut = "off";
defparam \Add0~117 .lut_mask = 64'h000000000000FF00;
defparam \Add0~117 .shared_arith = "off";

cyclonev_lcell_comb \internal_counter~8 (
	.dataa(!\always0~0_combout ),
	.datab(!\period_l_register[0]~q ),
	.datac(!\Add0~117_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\internal_counter~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \internal_counter~8 .extended_lut = "off";
defparam \internal_counter~8 .lut_mask = 64'hB1B1B1B1B1B1B1B1;
defparam \internal_counter~8 .shared_arith = "off";

cyclonev_lcell_comb \force_reload~0 (
	.dataa(!A_mem_baddr_3),
	.datab(!A_mem_baddr_4),
	.datac(!\period_l_wr_strobe~1_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\force_reload~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \force_reload~0 .extended_lut = "off";
defparam \force_reload~0 .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \force_reload~0 .shared_arith = "off";

dffeas force_reload(
	.clk(clk),
	.d(\force_reload~0_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\force_reload~q ),
	.prn(vcc));
defparam force_reload.is_wysiwyg = "true";
defparam force_reload.power_up = "low";

cyclonev_lcell_comb \Equal6~0 (
	.dataa(!A_mem_baddr_3),
	.datab(!A_mem_baddr_2),
	.datac(!A_mem_baddr_4),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal6~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal6~0 .extended_lut = "off";
defparam \Equal6~0 .lut_mask = 64'hFBFBFBFBFBFBFBFB;
defparam \Equal6~0 .shared_arith = "off";

cyclonev_lcell_comb control_wr_strobe(
	.dataa(!clr_break_line),
	.datab(!Equal2),
	.datac(!mem_used_1),
	.datad(!wait_latency_counter_1),
	.datae(!\period_l_wr_strobe~0_combout ),
	.dataf(!\Equal6~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\control_wr_strobe~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam control_wr_strobe.extended_lut = "off";
defparam control_wr_strobe.lut_mask = 64'hFFF7FFFFFFFFFFFF;
defparam control_wr_strobe.shared_arith = "off";

dffeas \control_register[1] (
	.clk(clk),
	.d(writedata[1]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\control_wr_strobe~combout ),
	.q(\control_register[1]~q ),
	.prn(vcc));
defparam \control_register[1] .is_wysiwyg = "true";
defparam \control_register[1] .power_up = "low";

cyclonev_lcell_comb \counter_is_running~0 (
	.dataa(!\force_reload~q ),
	.datab(!\counter_is_running~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\counter_is_running~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \counter_is_running~0 .extended_lut = "off";
defparam \counter_is_running~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \counter_is_running~0 .shared_arith = "off";

cyclonev_lcell_comb \counter_is_running~1 (
	.dataa(!writedata[2]),
	.datab(!writedata[3]),
	.datac(!\Equal0~6_combout ),
	.datad(!\control_wr_strobe~combout ),
	.datae(!\control_register[1]~q ),
	.dataf(!\counter_is_running~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\counter_is_running~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \counter_is_running~1 .extended_lut = "off";
defparam \counter_is_running~1 .lut_mask = 64'hDDF5FFFFFFFFFFFF;
defparam \counter_is_running~1 .shared_arith = "off";

dffeas counter_is_running(
	.clk(clk),
	.d(\counter_is_running~1_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\counter_is_running~q ),
	.prn(vcc));
defparam counter_is_running.is_wysiwyg = "true";
defparam counter_is_running.power_up = "low";

cyclonev_lcell_comb \always0~1 (
	.dataa(!\force_reload~q ),
	.datab(!\counter_is_running~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~1 .extended_lut = "off";
defparam \always0~1 .lut_mask = 64'h7777777777777777;
defparam \always0~1 .shared_arith = "off";

dffeas \internal_counter[0] (
	.clk(clk),
	.d(\internal_counter~8_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\internal_counter[0]~q ),
	.prn(vcc));
defparam \internal_counter[0] .is_wysiwyg = "true";
defparam \internal_counter[0] .power_up = "low";

cyclonev_lcell_comb \Add0~113 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\internal_counter[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~118 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~113_sumout ),
	.cout(\Add0~114 ),
	.shareout());
defparam \Add0~113 .extended_lut = "off";
defparam \Add0~113 .lut_mask = 64'h000000000000FF00;
defparam \Add0~113 .shared_arith = "off";

cyclonev_lcell_comb \internal_counter~7 (
	.dataa(!\always0~0_combout ),
	.datab(!\period_l_register[1]~q ),
	.datac(!\Add0~113_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\internal_counter~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \internal_counter~7 .extended_lut = "off";
defparam \internal_counter~7 .lut_mask = 64'hB1B1B1B1B1B1B1B1;
defparam \internal_counter~7 .shared_arith = "off";

dffeas \internal_counter[1] (
	.clk(clk),
	.d(\internal_counter~7_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\internal_counter[1]~q ),
	.prn(vcc));
defparam \internal_counter[1] .is_wysiwyg = "true";
defparam \internal_counter[1] .power_up = "low";

cyclonev_lcell_comb \Add0~109 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\internal_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~114 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~109_sumout ),
	.cout(\Add0~110 ),
	.shareout());
defparam \Add0~109 .extended_lut = "off";
defparam \Add0~109 .lut_mask = 64'h000000000000FF00;
defparam \Add0~109 .shared_arith = "off";

cyclonev_lcell_comb \internal_counter~6 (
	.dataa(!\always0~0_combout ),
	.datab(!\period_l_register[2]~q ),
	.datac(!\Add0~109_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\internal_counter~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \internal_counter~6 .extended_lut = "off";
defparam \internal_counter~6 .lut_mask = 64'hB1B1B1B1B1B1B1B1;
defparam \internal_counter~6 .shared_arith = "off";

dffeas \internal_counter[2] (
	.clk(clk),
	.d(\internal_counter~6_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\internal_counter[2]~q ),
	.prn(vcc));
defparam \internal_counter[2] .is_wysiwyg = "true";
defparam \internal_counter[2] .power_up = "low";

cyclonev_lcell_comb \Add0~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\internal_counter[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~110 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~57_sumout ),
	.cout(\Add0~58 ),
	.shareout());
defparam \Add0~57 .extended_lut = "off";
defparam \Add0~57 .lut_mask = 64'h000000000000FF00;
defparam \Add0~57 .shared_arith = "off";

cyclonev_lcell_comb \internal_counter~0 (
	.dataa(!\always0~0_combout ),
	.datab(!\period_l_register[3]~q ),
	.datac(!\Add0~57_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\internal_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \internal_counter~0 .extended_lut = "off";
defparam \internal_counter~0 .lut_mask = 64'hB1B1B1B1B1B1B1B1;
defparam \internal_counter~0 .shared_arith = "off";

dffeas \internal_counter[3] (
	.clk(clk),
	.d(\internal_counter~0_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\internal_counter[3]~q ),
	.prn(vcc));
defparam \internal_counter[3] .is_wysiwyg = "true";
defparam \internal_counter[3] .power_up = "low";

cyclonev_lcell_comb \Add0~125 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\internal_counter[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~125_sumout ),
	.cout(\Add0~126 ),
	.shareout());
defparam \Add0~125 .extended_lut = "off";
defparam \Add0~125 .lut_mask = 64'h00000000000000FF;
defparam \Add0~125 .shared_arith = "off";

dffeas \period_l_register[4] (
	.clk(clk),
	.d(writedata[4]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_l_wr_strobe~combout ),
	.q(\period_l_register[4]~q ),
	.prn(vcc));
defparam \period_l_register[4] .is_wysiwyg = "true";
defparam \period_l_register[4] .power_up = "low";

dffeas \internal_counter[4] (
	.clk(clk),
	.d(\Add0~125_sumout ),
	.asdata(\period_l_register[4]~q ),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always0~0_combout ),
	.ena(\always0~1_combout ),
	.q(\internal_counter[4]~q ),
	.prn(vcc));
defparam \internal_counter[4] .is_wysiwyg = "true";
defparam \internal_counter[4] .power_up = "low";

cyclonev_lcell_comb \Add0~121 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\internal_counter[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~126 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~121_sumout ),
	.cout(\Add0~122 ),
	.shareout());
defparam \Add0~121 .extended_lut = "off";
defparam \Add0~121 .lut_mask = 64'h00000000000000FF;
defparam \Add0~121 .shared_arith = "off";

dffeas \period_l_register[5] (
	.clk(clk),
	.d(writedata[5]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_l_wr_strobe~combout ),
	.q(\period_l_register[5]~q ),
	.prn(vcc));
defparam \period_l_register[5] .is_wysiwyg = "true";
defparam \period_l_register[5] .power_up = "low";

dffeas \internal_counter[5] (
	.clk(clk),
	.d(\Add0~121_sumout ),
	.asdata(\period_l_register[5]~q ),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always0~0_combout ),
	.ena(\always0~1_combout ),
	.q(\internal_counter[5]~q ),
	.prn(vcc));
defparam \internal_counter[5] .is_wysiwyg = "true";
defparam \internal_counter[5] .power_up = "low";

cyclonev_lcell_comb \Add0~105 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\internal_counter[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~122 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~105_sumout ),
	.cout(\Add0~106 ),
	.shareout());
defparam \Add0~105 .extended_lut = "off";
defparam \Add0~105 .lut_mask = 64'h000000000000FF00;
defparam \Add0~105 .shared_arith = "off";

cyclonev_lcell_comb \internal_counter~5 (
	.dataa(!\always0~0_combout ),
	.datab(!\period_l_register[6]~q ),
	.datac(!\Add0~105_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\internal_counter~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \internal_counter~5 .extended_lut = "off";
defparam \internal_counter~5 .lut_mask = 64'hB1B1B1B1B1B1B1B1;
defparam \internal_counter~5 .shared_arith = "off";

dffeas \internal_counter[6] (
	.clk(clk),
	.d(\internal_counter~5_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\internal_counter[6]~q ),
	.prn(vcc));
defparam \internal_counter[6] .is_wysiwyg = "true";
defparam \internal_counter[6] .power_up = "low";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\internal_counter[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~106 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h00000000000000FF;
defparam \Add0~5 .shared_arith = "off";

dffeas \period_l_register[7] (
	.clk(clk),
	.d(writedata[7]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_l_wr_strobe~combout ),
	.q(\period_l_register[7]~q ),
	.prn(vcc));
defparam \period_l_register[7] .is_wysiwyg = "true";
defparam \period_l_register[7] .power_up = "low";

dffeas \internal_counter[7] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(\period_l_register[7]~q ),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always0~0_combout ),
	.ena(\always0~1_combout ),
	.q(\internal_counter[7]~q ),
	.prn(vcc));
defparam \internal_counter[7] .is_wysiwyg = "true";
defparam \internal_counter[7] .power_up = "low";

cyclonev_lcell_comb \period_l_register[15]~1 (
	.dataa(!writedata[15]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\period_l_register[15]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \period_l_register[15]~1 .extended_lut = "off";
defparam \period_l_register[15]~1 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \period_l_register[15]~1 .shared_arith = "off";

dffeas \period_l_register[15] (
	.clk(clk),
	.d(\period_l_register[15]~1_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_l_wr_strobe~combout ),
	.q(\period_l_register[15]~q ),
	.prn(vcc));
defparam \period_l_register[15] .is_wysiwyg = "true";
defparam \period_l_register[15] .power_up = "low";

cyclonev_lcell_comb \period_l_register[14]~2 (
	.dataa(!writedata[14]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\period_l_register[14]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \period_l_register[14]~2 .extended_lut = "off";
defparam \period_l_register[14]~2 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \period_l_register[14]~2 .shared_arith = "off";

dffeas \period_l_register[14] (
	.clk(clk),
	.d(\period_l_register[14]~2_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_l_wr_strobe~combout ),
	.q(\period_l_register[14]~q ),
	.prn(vcc));
defparam \period_l_register[14] .is_wysiwyg = "true";
defparam \period_l_register[14] .power_up = "low";

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\internal_counter[10]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~98 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(\Add0~2 ),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h00000000000000FF;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\internal_counter[11]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout());
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h00000000000000FF;
defparam \Add0~29 .shared_arith = "off";

dffeas \period_l_register[11] (
	.clk(clk),
	.d(writedata[11]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_l_wr_strobe~combout ),
	.q(\period_l_register[11]~q ),
	.prn(vcc));
defparam \period_l_register[11] .is_wysiwyg = "true";
defparam \period_l_register[11] .power_up = "low";

dffeas \internal_counter[11] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(\period_l_register[11]~q ),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always0~0_combout ),
	.ena(\always0~1_combout ),
	.q(\internal_counter[11]~q ),
	.prn(vcc));
defparam \internal_counter[11] .is_wysiwyg = "true";
defparam \internal_counter[11] .power_up = "low";

cyclonev_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\internal_counter[12]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h00000000000000FF;
defparam \Add0~25 .shared_arith = "off";

dffeas \period_l_register[12] (
	.clk(clk),
	.d(writedata[12]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_l_wr_strobe~combout ),
	.q(\period_l_register[12]~q ),
	.prn(vcc));
defparam \period_l_register[12] .is_wysiwyg = "true";
defparam \period_l_register[12] .power_up = "low";

dffeas \internal_counter[12] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(\period_l_register[12]~q ),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always0~0_combout ),
	.ena(\always0~1_combout ),
	.q(\internal_counter[12]~q ),
	.prn(vcc));
defparam \internal_counter[12] .is_wysiwyg = "true";
defparam \internal_counter[12] .power_up = "low";

cyclonev_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\internal_counter[13]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h00000000000000FF;
defparam \Add0~21 .shared_arith = "off";

dffeas \period_l_register[13] (
	.clk(clk),
	.d(writedata[13]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_l_wr_strobe~combout ),
	.q(\period_l_register[13]~q ),
	.prn(vcc));
defparam \period_l_register[13] .is_wysiwyg = "true";
defparam \period_l_register[13] .power_up = "low";

dffeas \internal_counter[13] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(\period_l_register[13]~q ),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always0~0_combout ),
	.ena(\always0~1_combout ),
	.q(\internal_counter[13]~q ),
	.prn(vcc));
defparam \internal_counter[13] .is_wysiwyg = "true";
defparam \internal_counter[13] .power_up = "low";

cyclonev_lcell_comb \Add0~93 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\internal_counter[14]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~93_sumout ),
	.cout(\Add0~94 ),
	.shareout());
defparam \Add0~93 .extended_lut = "off";
defparam \Add0~93 .lut_mask = 64'h000000000000FF00;
defparam \Add0~93 .shared_arith = "off";

cyclonev_lcell_comb \internal_counter~2 (
	.dataa(!\always0~0_combout ),
	.datab(!\period_l_register[14]~q ),
	.datac(!\Add0~93_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\internal_counter~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \internal_counter~2 .extended_lut = "off";
defparam \internal_counter~2 .lut_mask = 64'hB1B1B1B1B1B1B1B1;
defparam \internal_counter~2 .shared_arith = "off";

dffeas \internal_counter[14] (
	.clk(clk),
	.d(\internal_counter~2_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\internal_counter[14]~q ),
	.prn(vcc));
defparam \internal_counter[14] .is_wysiwyg = "true";
defparam \internal_counter[14] .power_up = "low";

cyclonev_lcell_comb \Add0~89 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\internal_counter[15]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~94 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~89_sumout ),
	.cout(\Add0~90 ),
	.shareout());
defparam \Add0~89 .extended_lut = "off";
defparam \Add0~89 .lut_mask = 64'h000000000000FF00;
defparam \Add0~89 .shared_arith = "off";

cyclonev_lcell_comb \internal_counter~1 (
	.dataa(!\always0~0_combout ),
	.datab(!\period_l_register[15]~q ),
	.datac(!\Add0~89_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\internal_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \internal_counter~1 .extended_lut = "off";
defparam \internal_counter~1 .lut_mask = 64'hB1B1B1B1B1B1B1B1;
defparam \internal_counter~1 .shared_arith = "off";

dffeas \internal_counter[15] (
	.clk(clk),
	.d(\internal_counter~1_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\internal_counter[15]~q ),
	.prn(vcc));
defparam \internal_counter[15] .is_wysiwyg = "true";
defparam \internal_counter[15] .power_up = "low";

cyclonev_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\internal_counter[16]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~90 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h00000000000000FF;
defparam \Add0~17 .shared_arith = "off";

cyclonev_lcell_comb \Equal6~1 (
	.dataa(!A_mem_baddr_3),
	.datab(!A_mem_baddr_2),
	.datac(!A_mem_baddr_4),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal6~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal6~1 .extended_lut = "off";
defparam \Equal6~1 .lut_mask = 64'hF7F7F7F7F7F7F7F7;
defparam \Equal6~1 .shared_arith = "off";

cyclonev_lcell_comb period_h_wr_strobe(
	.dataa(!clr_break_line),
	.datab(!Equal2),
	.datac(!mem_used_1),
	.datad(!wait_latency_counter_1),
	.datae(!\period_l_wr_strobe~0_combout ),
	.dataf(!\Equal6~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\period_h_wr_strobe~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam period_h_wr_strobe.extended_lut = "off";
defparam period_h_wr_strobe.lut_mask = 64'hFFF7FFFFFFFFFFFF;
defparam period_h_wr_strobe.shared_arith = "off";

dffeas \period_h_register[0] (
	.clk(clk),
	.d(writedata[0]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_h_wr_strobe~combout ),
	.q(\period_h_register[0]~q ),
	.prn(vcc));
defparam \period_h_register[0] .is_wysiwyg = "true";
defparam \period_h_register[0] .power_up = "low";

dffeas \internal_counter[16] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(\period_h_register[0]~q ),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always0~0_combout ),
	.ena(\always0~1_combout ),
	.q(\internal_counter[16]~q ),
	.prn(vcc));
defparam \internal_counter[16] .is_wysiwyg = "true";
defparam \internal_counter[16] .power_up = "low";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\internal_counter[17]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h00000000000000FF;
defparam \Add0~13 .shared_arith = "off";

dffeas \period_h_register[1] (
	.clk(clk),
	.d(writedata[1]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_h_wr_strobe~combout ),
	.q(\period_h_register[1]~q ),
	.prn(vcc));
defparam \period_h_register[1] .is_wysiwyg = "true";
defparam \period_h_register[1] .power_up = "low";

dffeas \internal_counter[17] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(\period_h_register[1]~q ),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always0~0_combout ),
	.ena(\always0~1_combout ),
	.q(\internal_counter[17]~q ),
	.prn(vcc));
defparam \internal_counter[17] .is_wysiwyg = "true";
defparam \internal_counter[17] .power_up = "low";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\internal_counter[18]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h00000000000000FF;
defparam \Add0~9 .shared_arith = "off";

dffeas \period_h_register[2] (
	.clk(clk),
	.d(writedata[2]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_h_wr_strobe~combout ),
	.q(\period_h_register[2]~q ),
	.prn(vcc));
defparam \period_h_register[2] .is_wysiwyg = "true";
defparam \period_h_register[2] .power_up = "low";

dffeas \internal_counter[18] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(\period_h_register[2]~q ),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always0~0_combout ),
	.ena(\always0~1_combout ),
	.q(\internal_counter[18]~q ),
	.prn(vcc));
defparam \internal_counter[18] .is_wysiwyg = "true";
defparam \internal_counter[18] .power_up = "low";

cyclonev_lcell_comb \Equal0~0 (
	.dataa(!\internal_counter[18]~q ),
	.datab(!\internal_counter[17]~q ),
	.datac(!\internal_counter[16]~q ),
	.datad(!\internal_counter[13]~q ),
	.datae(!\internal_counter[12]~q ),
	.dataf(!\internal_counter[11]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~0 .extended_lut = "off";
defparam \Equal0~0 .lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam \Equal0~0 .shared_arith = "off";

cyclonev_lcell_comb \Add0~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\internal_counter[19]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~53_sumout ),
	.cout(\Add0~54 ),
	.shareout());
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h00000000000000FF;
defparam \Add0~53 .shared_arith = "off";

dffeas \period_h_register[3] (
	.clk(clk),
	.d(writedata[3]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_h_wr_strobe~combout ),
	.q(\period_h_register[3]~q ),
	.prn(vcc));
defparam \period_h_register[3] .is_wysiwyg = "true";
defparam \period_h_register[3] .power_up = "low";

dffeas \internal_counter[19] (
	.clk(clk),
	.d(\Add0~53_sumout ),
	.asdata(\period_h_register[3]~q ),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always0~0_combout ),
	.ena(\always0~1_combout ),
	.q(\internal_counter[19]~q ),
	.prn(vcc));
defparam \internal_counter[19] .is_wysiwyg = "true";
defparam \internal_counter[19] .power_up = "low";

cyclonev_lcell_comb \Add0~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\internal_counter[20]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~61_sumout ),
	.cout(\Add0~62 ),
	.shareout());
defparam \Add0~61 .extended_lut = "off";
defparam \Add0~61 .lut_mask = 64'h00000000000000FF;
defparam \Add0~61 .shared_arith = "off";

dffeas \period_h_register[4] (
	.clk(clk),
	.d(writedata[4]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_h_wr_strobe~combout ),
	.q(\period_h_register[4]~q ),
	.prn(vcc));
defparam \period_h_register[4] .is_wysiwyg = "true";
defparam \period_h_register[4] .power_up = "low";

dffeas \internal_counter[20] (
	.clk(clk),
	.d(\Add0~61_sumout ),
	.asdata(\period_h_register[4]~q ),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always0~0_combout ),
	.ena(\always0~1_combout ),
	.q(\internal_counter[20]~q ),
	.prn(vcc));
defparam \internal_counter[20] .is_wysiwyg = "true";
defparam \internal_counter[20] .power_up = "low";

cyclonev_lcell_comb \Add0~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\internal_counter[21]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~49_sumout ),
	.cout(\Add0~50 ),
	.shareout());
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h00000000000000FF;
defparam \Add0~49 .shared_arith = "off";

dffeas \period_h_register[5] (
	.clk(clk),
	.d(writedata[5]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_h_wr_strobe~combout ),
	.q(\period_h_register[5]~q ),
	.prn(vcc));
defparam \period_h_register[5] .is_wysiwyg = "true";
defparam \period_h_register[5] .power_up = "low";

dffeas \internal_counter[21] (
	.clk(clk),
	.d(\Add0~49_sumout ),
	.asdata(\period_h_register[5]~q ),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always0~0_combout ),
	.ena(\always0~1_combout ),
	.q(\internal_counter[21]~q ),
	.prn(vcc));
defparam \internal_counter[21] .is_wysiwyg = "true";
defparam \internal_counter[21] .power_up = "low";

cyclonev_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\internal_counter[22]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout());
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h00000000000000FF;
defparam \Add0~45 .shared_arith = "off";

dffeas \period_h_register[6] (
	.clk(clk),
	.d(writedata[6]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_h_wr_strobe~combout ),
	.q(\period_h_register[6]~q ),
	.prn(vcc));
defparam \period_h_register[6] .is_wysiwyg = "true";
defparam \period_h_register[6] .power_up = "low";

dffeas \internal_counter[22] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(\period_h_register[6]~q ),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always0~0_combout ),
	.ena(\always0~1_combout ),
	.q(\internal_counter[22]~q ),
	.prn(vcc));
defparam \internal_counter[22] .is_wysiwyg = "true";
defparam \internal_counter[22] .power_up = "low";

cyclonev_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\internal_counter[23]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout());
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h00000000000000FF;
defparam \Add0~41 .shared_arith = "off";

dffeas \period_h_register[7] (
	.clk(clk),
	.d(writedata[7]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_h_wr_strobe~combout ),
	.q(\period_h_register[7]~q ),
	.prn(vcc));
defparam \period_h_register[7] .is_wysiwyg = "true";
defparam \period_h_register[7] .power_up = "low";

dffeas \internal_counter[23] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(\period_h_register[7]~q ),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always0~0_combout ),
	.ena(\always0~1_combout ),
	.q(\internal_counter[23]~q ),
	.prn(vcc));
defparam \internal_counter[23] .is_wysiwyg = "true";
defparam \internal_counter[23] .power_up = "low";

cyclonev_lcell_comb \Add0~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\internal_counter[24]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~69_sumout ),
	.cout(\Add0~70 ),
	.shareout());
defparam \Add0~69 .extended_lut = "off";
defparam \Add0~69 .lut_mask = 64'h00000000000000FF;
defparam \Add0~69 .shared_arith = "off";

dffeas \period_h_register[8] (
	.clk(clk),
	.d(writedata[8]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_h_wr_strobe~combout ),
	.q(\period_h_register[8]~q ),
	.prn(vcc));
defparam \period_h_register[8] .is_wysiwyg = "true";
defparam \period_h_register[8] .power_up = "low";

dffeas \internal_counter[24] (
	.clk(clk),
	.d(\Add0~69_sumout ),
	.asdata(\period_h_register[8]~q ),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always0~0_combout ),
	.ena(\always0~1_combout ),
	.q(\internal_counter[24]~q ),
	.prn(vcc));
defparam \internal_counter[24] .is_wysiwyg = "true";
defparam \internal_counter[24] .power_up = "low";

cyclonev_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\internal_counter[25]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~70 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout());
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h00000000000000FF;
defparam \Add0~37 .shared_arith = "off";

dffeas \period_h_register[9] (
	.clk(clk),
	.d(writedata[9]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_h_wr_strobe~combout ),
	.q(\period_h_register[9]~q ),
	.prn(vcc));
defparam \period_h_register[9] .is_wysiwyg = "true";
defparam \period_h_register[9] .power_up = "low";

dffeas \internal_counter[25] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(\period_h_register[9]~q ),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always0~0_combout ),
	.ena(\always0~1_combout ),
	.q(\internal_counter[25]~q ),
	.prn(vcc));
defparam \internal_counter[25] .is_wysiwyg = "true";
defparam \internal_counter[25] .power_up = "low";

cyclonev_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\internal_counter[26]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout());
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h00000000000000FF;
defparam \Add0~33 .shared_arith = "off";

dffeas \period_h_register[10] (
	.clk(clk),
	.d(writedata[10]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_h_wr_strobe~combout ),
	.q(\period_h_register[10]~q ),
	.prn(vcc));
defparam \period_h_register[10] .is_wysiwyg = "true";
defparam \period_h_register[10] .power_up = "low";

dffeas \internal_counter[26] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(\period_h_register[10]~q ),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always0~0_combout ),
	.ena(\always0~1_combout ),
	.q(\internal_counter[26]~q ),
	.prn(vcc));
defparam \internal_counter[26] .is_wysiwyg = "true";
defparam \internal_counter[26] .power_up = "low";

cyclonev_lcell_comb \Equal0~1 (
	.dataa(!\internal_counter[26]~q ),
	.datab(!\internal_counter[25]~q ),
	.datac(!\internal_counter[23]~q ),
	.datad(!\internal_counter[22]~q ),
	.datae(!\internal_counter[21]~q ),
	.dataf(!\internal_counter[19]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~1 .extended_lut = "off";
defparam \Equal0~1 .lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam \Equal0~1 .shared_arith = "off";

cyclonev_lcell_comb \Add0~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\internal_counter[27]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~65_sumout ),
	.cout(\Add0~66 ),
	.shareout());
defparam \Add0~65 .extended_lut = "off";
defparam \Add0~65 .lut_mask = 64'h00000000000000FF;
defparam \Add0~65 .shared_arith = "off";

dffeas \period_h_register[11] (
	.clk(clk),
	.d(writedata[11]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_h_wr_strobe~combout ),
	.q(\period_h_register[11]~q ),
	.prn(vcc));
defparam \period_h_register[11] .is_wysiwyg = "true";
defparam \period_h_register[11] .power_up = "low";

dffeas \internal_counter[27] (
	.clk(clk),
	.d(\Add0~65_sumout ),
	.asdata(\period_h_register[11]~q ),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always0~0_combout ),
	.ena(\always0~1_combout ),
	.q(\internal_counter[27]~q ),
	.prn(vcc));
defparam \internal_counter[27] .is_wysiwyg = "true";
defparam \internal_counter[27] .power_up = "low";

cyclonev_lcell_comb \Add0~85 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\internal_counter[28]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~66 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~85_sumout ),
	.cout(\Add0~86 ),
	.shareout());
defparam \Add0~85 .extended_lut = "off";
defparam \Add0~85 .lut_mask = 64'h00000000000000FF;
defparam \Add0~85 .shared_arith = "off";

dffeas \period_h_register[12] (
	.clk(clk),
	.d(writedata[12]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_h_wr_strobe~combout ),
	.q(\period_h_register[12]~q ),
	.prn(vcc));
defparam \period_h_register[12] .is_wysiwyg = "true";
defparam \period_h_register[12] .power_up = "low";

dffeas \internal_counter[28] (
	.clk(clk),
	.d(\Add0~85_sumout ),
	.asdata(\period_h_register[12]~q ),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always0~0_combout ),
	.ena(\always0~1_combout ),
	.q(\internal_counter[28]~q ),
	.prn(vcc));
defparam \internal_counter[28] .is_wysiwyg = "true";
defparam \internal_counter[28] .power_up = "low";

cyclonev_lcell_comb \Add0~81 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\internal_counter[29]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~86 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~81_sumout ),
	.cout(\Add0~82 ),
	.shareout());
defparam \Add0~81 .extended_lut = "off";
defparam \Add0~81 .lut_mask = 64'h00000000000000FF;
defparam \Add0~81 .shared_arith = "off";

dffeas \period_h_register[13] (
	.clk(clk),
	.d(writedata[13]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_h_wr_strobe~combout ),
	.q(\period_h_register[13]~q ),
	.prn(vcc));
defparam \period_h_register[13] .is_wysiwyg = "true";
defparam \period_h_register[13] .power_up = "low";

dffeas \internal_counter[29] (
	.clk(clk),
	.d(\Add0~81_sumout ),
	.asdata(\period_h_register[13]~q ),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always0~0_combout ),
	.ena(\always0~1_combout ),
	.q(\internal_counter[29]~q ),
	.prn(vcc));
defparam \internal_counter[29] .is_wysiwyg = "true";
defparam \internal_counter[29] .power_up = "low";

cyclonev_lcell_comb \Add0~77 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\internal_counter[30]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~82 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~77_sumout ),
	.cout(\Add0~78 ),
	.shareout());
defparam \Add0~77 .extended_lut = "off";
defparam \Add0~77 .lut_mask = 64'h00000000000000FF;
defparam \Add0~77 .shared_arith = "off";

dffeas \period_h_register[14] (
	.clk(clk),
	.d(writedata[14]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_h_wr_strobe~combout ),
	.q(\period_h_register[14]~q ),
	.prn(vcc));
defparam \period_h_register[14] .is_wysiwyg = "true";
defparam \period_h_register[14] .power_up = "low";

dffeas \internal_counter[30] (
	.clk(clk),
	.d(\Add0~77_sumout ),
	.asdata(\period_h_register[14]~q ),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always0~0_combout ),
	.ena(\always0~1_combout ),
	.q(\internal_counter[30]~q ),
	.prn(vcc));
defparam \internal_counter[30] .is_wysiwyg = "true";
defparam \internal_counter[30] .power_up = "low";

cyclonev_lcell_comb \Add0~73 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\internal_counter[31]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~78 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~73_sumout ),
	.cout(),
	.shareout());
defparam \Add0~73 .extended_lut = "off";
defparam \Add0~73 .lut_mask = 64'h00000000000000FF;
defparam \Add0~73 .shared_arith = "off";

dffeas \period_h_register[15] (
	.clk(clk),
	.d(writedata[15]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_h_wr_strobe~combout ),
	.q(\period_h_register[15]~q ),
	.prn(vcc));
defparam \period_h_register[15] .is_wysiwyg = "true";
defparam \period_h_register[15] .power_up = "low";

dffeas \internal_counter[31] (
	.clk(clk),
	.d(\Add0~73_sumout ),
	.asdata(\period_h_register[15]~q ),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always0~0_combout ),
	.ena(\always0~1_combout ),
	.q(\internal_counter[31]~q ),
	.prn(vcc));
defparam \internal_counter[31] .is_wysiwyg = "true";
defparam \internal_counter[31] .power_up = "low";

cyclonev_lcell_comb \Equal0~2 (
	.dataa(!\internal_counter[24]~q ),
	.datab(!\internal_counter[31]~q ),
	.datac(!\internal_counter[30]~q ),
	.datad(!\internal_counter[29]~q ),
	.datae(!\internal_counter[28]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~2 .extended_lut = "off";
defparam \Equal0~2 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \Equal0~2 .shared_arith = "off";

cyclonev_lcell_comb \period_l_register[8]~4 (
	.dataa(!writedata[8]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\period_l_register[8]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \period_l_register[8]~4 .extended_lut = "off";
defparam \period_l_register[8]~4 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \period_l_register[8]~4 .shared_arith = "off";

dffeas \period_l_register[8] (
	.clk(clk),
	.d(\period_l_register[8]~4_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_l_wr_strobe~combout ),
	.q(\period_l_register[8]~q ),
	.prn(vcc));
defparam \period_l_register[8] .is_wysiwyg = "true";
defparam \period_l_register[8] .power_up = "low";

cyclonev_lcell_comb \Add0~101 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\internal_counter[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~101_sumout ),
	.cout(\Add0~102 ),
	.shareout());
defparam \Add0~101 .extended_lut = "off";
defparam \Add0~101 .lut_mask = 64'h000000000000FF00;
defparam \Add0~101 .shared_arith = "off";

cyclonev_lcell_comb \internal_counter~4 (
	.dataa(!\always0~0_combout ),
	.datab(!\period_l_register[8]~q ),
	.datac(!\Add0~101_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\internal_counter~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \internal_counter~4 .extended_lut = "off";
defparam \internal_counter~4 .lut_mask = 64'hB1B1B1B1B1B1B1B1;
defparam \internal_counter~4 .shared_arith = "off";

dffeas \internal_counter[8] (
	.clk(clk),
	.d(\internal_counter~4_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\internal_counter[8]~q ),
	.prn(vcc));
defparam \internal_counter[8] .is_wysiwyg = "true";
defparam \internal_counter[8] .power_up = "low";

cyclonev_lcell_comb \Equal0~3 (
	.dataa(!\internal_counter[15]~q ),
	.datab(!\internal_counter[14]~q ),
	.datac(!\internal_counter[9]~q ),
	.datad(!\internal_counter[8]~q ),
	.datae(!\internal_counter[6]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~3 .extended_lut = "off";
defparam \Equal0~3 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \Equal0~3 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~4 (
	.dataa(!\internal_counter[2]~q ),
	.datab(!\internal_counter[1]~q ),
	.datac(!\internal_counter[0]~q ),
	.datad(!\internal_counter[5]~q ),
	.datae(!\internal_counter[4]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~4 .extended_lut = "off";
defparam \Equal0~4 .lut_mask = 64'hFFFFFF7FFFFFFF7F;
defparam \Equal0~4 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~5 (
	.dataa(!\internal_counter[3]~q ),
	.datab(!\internal_counter[20]~q ),
	.datac(!\internal_counter[27]~q ),
	.datad(!\Equal0~2_combout ),
	.datae(!\Equal0~3_combout ),
	.dataf(!\Equal0~4_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~5 .extended_lut = "off";
defparam \Equal0~5 .lut_mask = 64'hFDFFFFFFFFFFFFFF;
defparam \Equal0~5 .shared_arith = "off";

cyclonev_lcell_comb \always0~0 (
	.dataa(!\internal_counter[10]~q ),
	.datab(!\internal_counter[7]~q ),
	.datac(!\Equal0~0_combout ),
	.datad(!\Equal0~1_combout ),
	.datae(!\Equal0~5_combout ),
	.dataf(!\force_reload~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'hEFFFFFFFFFFFFFFF;
defparam \always0~0 .shared_arith = "off";

cyclonev_lcell_comb \period_l_register[9]~3 (
	.dataa(!writedata[9]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\period_l_register[9]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \period_l_register[9]~3 .extended_lut = "off";
defparam \period_l_register[9]~3 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \period_l_register[9]~3 .shared_arith = "off";

dffeas \period_l_register[9] (
	.clk(clk),
	.d(\period_l_register[9]~3_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_l_wr_strobe~combout ),
	.q(\period_l_register[9]~q ),
	.prn(vcc));
defparam \period_l_register[9] .is_wysiwyg = "true";
defparam \period_l_register[9] .power_up = "low";

cyclonev_lcell_comb \Add0~97 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\internal_counter[9]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~102 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~97_sumout ),
	.cout(\Add0~98 ),
	.shareout());
defparam \Add0~97 .extended_lut = "off";
defparam \Add0~97 .lut_mask = 64'h000000000000FF00;
defparam \Add0~97 .shared_arith = "off";

cyclonev_lcell_comb \internal_counter~3 (
	.dataa(!\always0~0_combout ),
	.datab(!\period_l_register[9]~q ),
	.datac(!\Add0~97_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\internal_counter~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \internal_counter~3 .extended_lut = "off";
defparam \internal_counter~3 .lut_mask = 64'hB1B1B1B1B1B1B1B1;
defparam \internal_counter~3 .shared_arith = "off";

dffeas \internal_counter[9] (
	.clk(clk),
	.d(\internal_counter~3_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\internal_counter[9]~q ),
	.prn(vcc));
defparam \internal_counter[9] .is_wysiwyg = "true";
defparam \internal_counter[9] .power_up = "low";

dffeas \period_l_register[10] (
	.clk(clk),
	.d(writedata[10]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_l_wr_strobe~combout ),
	.q(\period_l_register[10]~q ),
	.prn(vcc));
defparam \period_l_register[10] .is_wysiwyg = "true";
defparam \period_l_register[10] .power_up = "low";

dffeas \internal_counter[10] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(\period_l_register[10]~q ),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always0~0_combout ),
	.ena(\always0~1_combout ),
	.q(\internal_counter[10]~q ),
	.prn(vcc));
defparam \internal_counter[10] .is_wysiwyg = "true";
defparam \internal_counter[10] .power_up = "low";

cyclonev_lcell_comb \Equal0~6 (
	.dataa(!\internal_counter[10]~q ),
	.datab(!\internal_counter[7]~q ),
	.datac(!\Equal0~0_combout ),
	.datad(!\Equal0~1_combout ),
	.datae(!\Equal0~5_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~6 .extended_lut = "off";
defparam \Equal0~6 .lut_mask = 64'hEFFFFFFFEFFFFFFF;
defparam \Equal0~6 .shared_arith = "off";

dffeas delayed_unxcounter_is_zeroxx0(
	.clk(clk),
	.d(\Equal0~6_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delayed_unxcounter_is_zeroxx0~q ),
	.prn(vcc));
defparam delayed_unxcounter_is_zeroxx0.is_wysiwyg = "true";
defparam delayed_unxcounter_is_zeroxx0.power_up = "low";

cyclonev_lcell_comb \timeout_occurred~0 (
	.dataa(!timeout_occurred1),
	.datab(!\status_wr_strobe~0_combout ),
	.datac(!\delayed_unxcounter_is_zeroxx0~q ),
	.datad(!\Equal0~6_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\timeout_occurred~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \timeout_occurred~0 .extended_lut = "off";
defparam \timeout_occurred~0 .lut_mask = 64'hFDFFFDFFFDFFFDFF;
defparam \timeout_occurred~0 .shared_arith = "off";

cyclonev_lcell_comb \counter_snapshot[0]~0 (
	.dataa(!\internal_counter[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\counter_snapshot[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \counter_snapshot[0]~0 .extended_lut = "off";
defparam \counter_snapshot[0]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \counter_snapshot[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal6~3 (
	.dataa(!A_mem_baddr_3),
	.datab(!A_mem_baddr_4),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal6~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal6~3 .extended_lut = "off";
defparam \Equal6~3 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \Equal6~3 .shared_arith = "off";

cyclonev_lcell_comb \snap_strobe~0 (
	.dataa(!clr_break_line),
	.datab(!Equal2),
	.datac(!mem_used_1),
	.datad(!wait_latency_counter_1),
	.datae(!\period_l_wr_strobe~0_combout ),
	.dataf(!\Equal6~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\snap_strobe~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \snap_strobe~0 .extended_lut = "off";
defparam \snap_strobe~0 .lut_mask = 64'hFFF7FFFFFFFFFFFF;
defparam \snap_strobe~0 .shared_arith = "off";

dffeas \counter_snapshot[0] (
	.clk(clk),
	.d(\counter_snapshot[0]~0_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[0]~q ),
	.prn(vcc));
defparam \counter_snapshot[0] .is_wysiwyg = "true";
defparam \counter_snapshot[0] .power_up = "low";

cyclonev_lcell_comb \Equal6~4 (
	.dataa(!A_mem_baddr_2),
	.datab(!\Equal6~3_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal6~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal6~4 .extended_lut = "off";
defparam \Equal6~4 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \Equal6~4 .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[0]~0 (
	.dataa(!\period_l_register[0]~q ),
	.datab(!\Equal6~2_combout ),
	.datac(!\counter_snapshot[0]~q ),
	.datad(!\Equal6~4_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[0]~0 .extended_lut = "off";
defparam \read_mux_out[0]~0 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \read_mux_out[0]~0 .shared_arith = "off";

dffeas \counter_snapshot[16] (
	.clk(clk),
	.d(\internal_counter[16]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[16]~q ),
	.prn(vcc));
defparam \counter_snapshot[16] .is_wysiwyg = "true";
defparam \counter_snapshot[16] .power_up = "low";

cyclonev_lcell_comb \read_mux_out[0]~1 (
	.dataa(!A_mem_baddr_3),
	.datab(!A_mem_baddr_2),
	.datac(!A_mem_baddr_4),
	.datad(!timeout_occurred1),
	.datae(!control_register_0),
	.dataf(!\counter_snapshot[16]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[0]~1 .extended_lut = "off";
defparam \read_mux_out[0]~1 .lut_mask = 64'hBEFFFFFFFFFFFFFF;
defparam \read_mux_out[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[0] (
	.dataa(!\period_h_register[0]~q ),
	.datab(!\Equal6~1_combout ),
	.datac(!\read_mux_out[0]~0_combout ),
	.datad(!\read_mux_out[0]~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[0]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[0] .extended_lut = "off";
defparam \read_mux_out[0] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \read_mux_out[0] .shared_arith = "off";

cyclonev_lcell_comb \counter_snapshot[1]~1 (
	.dataa(!\internal_counter[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\counter_snapshot[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \counter_snapshot[1]~1 .extended_lut = "off";
defparam \counter_snapshot[1]~1 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \counter_snapshot[1]~1 .shared_arith = "off";

dffeas \counter_snapshot[1] (
	.clk(clk),
	.d(\counter_snapshot[1]~1_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[1]~q ),
	.prn(vcc));
defparam \counter_snapshot[1] .is_wysiwyg = "true";
defparam \counter_snapshot[1] .power_up = "low";

cyclonev_lcell_comb \read_mux_out[1]~2 (
	.dataa(!\period_l_register[1]~q ),
	.datab(!\Equal6~2_combout ),
	.datac(!\Equal6~4_combout ),
	.datad(!\counter_snapshot[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[1]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[1]~2 .extended_lut = "off";
defparam \read_mux_out[1]~2 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \read_mux_out[1]~2 .shared_arith = "off";

dffeas \counter_snapshot[17] (
	.clk(clk),
	.d(\internal_counter[17]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[17]~q ),
	.prn(vcc));
defparam \counter_snapshot[17] .is_wysiwyg = "true";
defparam \counter_snapshot[17] .power_up = "low";

cyclonev_lcell_comb \read_mux_out[1]~3 (
	.dataa(!A_mem_baddr_3),
	.datab(!A_mem_baddr_2),
	.datac(!A_mem_baddr_4),
	.datad(!\counter_is_running~q ),
	.datae(!\control_register[1]~q ),
	.dataf(!\counter_snapshot[17]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[1]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[1]~3 .extended_lut = "off";
defparam \read_mux_out[1]~3 .lut_mask = 64'hBEFFFFFFFFFFFFFF;
defparam \read_mux_out[1]~3 .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[1] (
	.dataa(!\period_h_register[1]~q ),
	.datab(!\Equal6~1_combout ),
	.datac(!\read_mux_out[1]~2_combout ),
	.datad(!\read_mux_out[1]~3_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[1]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[1] .extended_lut = "off";
defparam \read_mux_out[1] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \read_mux_out[1] .shared_arith = "off";

cyclonev_lcell_comb \counter_snapshot[2]~2 (
	.dataa(!\internal_counter[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\counter_snapshot[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \counter_snapshot[2]~2 .extended_lut = "off";
defparam \counter_snapshot[2]~2 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \counter_snapshot[2]~2 .shared_arith = "off";

dffeas \counter_snapshot[2] (
	.clk(clk),
	.d(\counter_snapshot[2]~2_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[2]~q ),
	.prn(vcc));
defparam \counter_snapshot[2] .is_wysiwyg = "true";
defparam \counter_snapshot[2] .power_up = "low";

cyclonev_lcell_comb \read_mux_out[2]~4 (
	.dataa(!\period_l_register[2]~q ),
	.datab(!\Equal6~2_combout ),
	.datac(!\Equal6~4_combout ),
	.datad(!\counter_snapshot[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[2]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[2]~4 .extended_lut = "off";
defparam \read_mux_out[2]~4 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \read_mux_out[2]~4 .shared_arith = "off";

cyclonev_lcell_comb \Equal6~5 (
	.dataa(!A_mem_baddr_2),
	.datab(!\Equal6~3_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal6~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal6~5 .extended_lut = "off";
defparam \Equal6~5 .lut_mask = 64'h7777777777777777;
defparam \Equal6~5 .shared_arith = "off";

dffeas \counter_snapshot[18] (
	.clk(clk),
	.d(\internal_counter[18]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[18]~q ),
	.prn(vcc));
defparam \counter_snapshot[18] .is_wysiwyg = "true";
defparam \counter_snapshot[18] .power_up = "low";

dffeas \control_register[2] (
	.clk(clk),
	.d(writedata[2]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\control_wr_strobe~combout ),
	.q(\control_register[2]~q ),
	.prn(vcc));
defparam \control_register[2] .is_wysiwyg = "true";
defparam \control_register[2] .power_up = "low";

cyclonev_lcell_comb \read_mux_out[2]~5 (
	.dataa(!\Equal6~0_combout ),
	.datab(!\Equal6~5_combout ),
	.datac(!\counter_snapshot[18]~q ),
	.datad(!\control_register[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[2]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[2]~5 .extended_lut = "off";
defparam \read_mux_out[2]~5 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \read_mux_out[2]~5 .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[2] (
	.dataa(!\period_h_register[2]~q ),
	.datab(!\Equal6~1_combout ),
	.datac(!\read_mux_out[2]~4_combout ),
	.datad(!\read_mux_out[2]~5_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[2]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[2] .extended_lut = "off";
defparam \read_mux_out[2] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \read_mux_out[2] .shared_arith = "off";

cyclonev_lcell_comb \counter_snapshot[3]~3 (
	.dataa(!\internal_counter[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\counter_snapshot[3]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \counter_snapshot[3]~3 .extended_lut = "off";
defparam \counter_snapshot[3]~3 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \counter_snapshot[3]~3 .shared_arith = "off";

dffeas \counter_snapshot[3] (
	.clk(clk),
	.d(\counter_snapshot[3]~3_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[3]~q ),
	.prn(vcc));
defparam \counter_snapshot[3] .is_wysiwyg = "true";
defparam \counter_snapshot[3] .power_up = "low";

cyclonev_lcell_comb \read_mux_out[3]~6 (
	.dataa(!\period_l_register[3]~q ),
	.datab(!\Equal6~2_combout ),
	.datac(!\Equal6~4_combout ),
	.datad(!\counter_snapshot[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[3]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[3]~6 .extended_lut = "off";
defparam \read_mux_out[3]~6 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \read_mux_out[3]~6 .shared_arith = "off";

dffeas \counter_snapshot[19] (
	.clk(clk),
	.d(\internal_counter[19]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[19]~q ),
	.prn(vcc));
defparam \counter_snapshot[19] .is_wysiwyg = "true";
defparam \counter_snapshot[19] .power_up = "low";

dffeas \control_register[3] (
	.clk(clk),
	.d(writedata[3]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\control_wr_strobe~combout ),
	.q(\control_register[3]~q ),
	.prn(vcc));
defparam \control_register[3] .is_wysiwyg = "true";
defparam \control_register[3] .power_up = "low";

cyclonev_lcell_comb \read_mux_out[3]~7 (
	.dataa(!\Equal6~0_combout ),
	.datab(!\Equal6~5_combout ),
	.datac(!\counter_snapshot[19]~q ),
	.datad(!\control_register[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[3]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[3]~7 .extended_lut = "off";
defparam \read_mux_out[3]~7 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \read_mux_out[3]~7 .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[3] (
	.dataa(!\period_h_register[3]~q ),
	.datab(!\Equal6~1_combout ),
	.datac(!\read_mux_out[3]~6_combout ),
	.datad(!\read_mux_out[3]~7_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[3]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[3] .extended_lut = "off";
defparam \read_mux_out[3] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \read_mux_out[3] .shared_arith = "off";

dffeas \counter_snapshot[4] (
	.clk(clk),
	.d(\internal_counter[4]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[4]~q ),
	.prn(vcc));
defparam \counter_snapshot[4] .is_wysiwyg = "true";
defparam \counter_snapshot[4] .power_up = "low";

dffeas \counter_snapshot[20] (
	.clk(clk),
	.d(\internal_counter[20]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[20]~q ),
	.prn(vcc));
defparam \counter_snapshot[20] .is_wysiwyg = "true";
defparam \counter_snapshot[20] .power_up = "low";

cyclonev_lcell_comb \read_mux_out[4]~52 (
	.dataa(!A_mem_baddr_2),
	.datab(!A_mem_baddr_3),
	.datac(!\counter_snapshot[4]~q ),
	.datad(!\counter_snapshot[20]~q ),
	.datae(!A_mem_baddr_4),
	.dataf(!\period_h_register[4]~q ),
	.datag(!\period_l_register[4]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[4]~52_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[4]~52 .extended_lut = "on";
defparam \read_mux_out[4]~52 .lut_mask = 64'hFFF6FFF6FFF6FFF6;
defparam \read_mux_out[4]~52 .shared_arith = "off";

dffeas \counter_snapshot[5] (
	.clk(clk),
	.d(\internal_counter[5]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[5]~q ),
	.prn(vcc));
defparam \counter_snapshot[5] .is_wysiwyg = "true";
defparam \counter_snapshot[5] .power_up = "low";

dffeas \counter_snapshot[21] (
	.clk(clk),
	.d(\internal_counter[21]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[21]~q ),
	.prn(vcc));
defparam \counter_snapshot[21] .is_wysiwyg = "true";
defparam \counter_snapshot[21] .power_up = "low";

cyclonev_lcell_comb \read_mux_out[5]~48 (
	.dataa(!A_mem_baddr_2),
	.datab(!A_mem_baddr_3),
	.datac(!\counter_snapshot[5]~q ),
	.datad(!\counter_snapshot[21]~q ),
	.datae(!A_mem_baddr_4),
	.dataf(!\period_h_register[5]~q ),
	.datag(!\period_l_register[5]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[5]~48_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[5]~48 .extended_lut = "on";
defparam \read_mux_out[5]~48 .lut_mask = 64'hFFF6FFF6FFF6FFF6;
defparam \read_mux_out[5]~48 .shared_arith = "off";

cyclonev_lcell_comb \counter_snapshot[6]~4 (
	.dataa(!\internal_counter[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\counter_snapshot[6]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \counter_snapshot[6]~4 .extended_lut = "off";
defparam \counter_snapshot[6]~4 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \counter_snapshot[6]~4 .shared_arith = "off";

dffeas \counter_snapshot[6] (
	.clk(clk),
	.d(\counter_snapshot[6]~4_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[6]~q ),
	.prn(vcc));
defparam \counter_snapshot[6] .is_wysiwyg = "true";
defparam \counter_snapshot[6] .power_up = "low";

dffeas \counter_snapshot[22] (
	.clk(clk),
	.d(\internal_counter[22]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[22]~q ),
	.prn(vcc));
defparam \counter_snapshot[22] .is_wysiwyg = "true";
defparam \counter_snapshot[22] .power_up = "low";

cyclonev_lcell_comb \read_mux_out[6]~44 (
	.dataa(!A_mem_baddr_2),
	.datab(!A_mem_baddr_3),
	.datac(!\counter_snapshot[6]~q ),
	.datad(!\counter_snapshot[22]~q ),
	.datae(!A_mem_baddr_4),
	.dataf(!\period_h_register[6]~q ),
	.datag(!\period_l_register[6]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[6]~44_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[6]~44 .extended_lut = "on";
defparam \read_mux_out[6]~44 .lut_mask = 64'hFF6FFFF6FF6FFFF6;
defparam \read_mux_out[6]~44 .shared_arith = "off";

dffeas \counter_snapshot[7] (
	.clk(clk),
	.d(\internal_counter[7]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[7]~q ),
	.prn(vcc));
defparam \counter_snapshot[7] .is_wysiwyg = "true";
defparam \counter_snapshot[7] .power_up = "low";

dffeas \counter_snapshot[23] (
	.clk(clk),
	.d(\internal_counter[23]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[23]~q ),
	.prn(vcc));
defparam \counter_snapshot[23] .is_wysiwyg = "true";
defparam \counter_snapshot[23] .power_up = "low";

cyclonev_lcell_comb \read_mux_out[7]~40 (
	.dataa(!A_mem_baddr_2),
	.datab(!A_mem_baddr_3),
	.datac(!\counter_snapshot[7]~q ),
	.datad(!\counter_snapshot[23]~q ),
	.datae(!A_mem_baddr_4),
	.dataf(!\period_h_register[7]~q ),
	.datag(!\period_l_register[7]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[7]~40_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[7]~40 .extended_lut = "on";
defparam \read_mux_out[7]~40 .lut_mask = 64'hFFF6FFF6FFF6FFF6;
defparam \read_mux_out[7]~40 .shared_arith = "off";

dffeas \counter_snapshot[11] (
	.clk(clk),
	.d(\internal_counter[11]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[11]~q ),
	.prn(vcc));
defparam \counter_snapshot[11] .is_wysiwyg = "true";
defparam \counter_snapshot[11] .power_up = "low";

dffeas \counter_snapshot[27] (
	.clk(clk),
	.d(\internal_counter[27]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[27]~q ),
	.prn(vcc));
defparam \counter_snapshot[27] .is_wysiwyg = "true";
defparam \counter_snapshot[27] .power_up = "low";

cyclonev_lcell_comb \read_mux_out[11]~36 (
	.dataa(!A_mem_baddr_2),
	.datab(!A_mem_baddr_3),
	.datac(!\counter_snapshot[11]~q ),
	.datad(!\counter_snapshot[27]~q ),
	.datae(!A_mem_baddr_4),
	.dataf(!\period_h_register[11]~q ),
	.datag(!\period_l_register[11]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[11]~36_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[11]~36 .extended_lut = "on";
defparam \read_mux_out[11]~36 .lut_mask = 64'hFFF6FFF6FFF6FFF6;
defparam \read_mux_out[11]~36 .shared_arith = "off";

dffeas \counter_snapshot[10] (
	.clk(clk),
	.d(\internal_counter[10]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[10]~q ),
	.prn(vcc));
defparam \counter_snapshot[10] .is_wysiwyg = "true";
defparam \counter_snapshot[10] .power_up = "low";

dffeas \counter_snapshot[26] (
	.clk(clk),
	.d(\internal_counter[26]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[26]~q ),
	.prn(vcc));
defparam \counter_snapshot[26] .is_wysiwyg = "true";
defparam \counter_snapshot[26] .power_up = "low";

cyclonev_lcell_comb \read_mux_out[10]~32 (
	.dataa(!A_mem_baddr_2),
	.datab(!A_mem_baddr_3),
	.datac(!\counter_snapshot[10]~q ),
	.datad(!\counter_snapshot[26]~q ),
	.datae(!A_mem_baddr_4),
	.dataf(!\period_h_register[10]~q ),
	.datag(!\period_l_register[10]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[10]~32_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[10]~32 .extended_lut = "on";
defparam \read_mux_out[10]~32 .lut_mask = 64'hFFF6FFF6FFF6FFF6;
defparam \read_mux_out[10]~32 .shared_arith = "off";

cyclonev_lcell_comb \counter_snapshot[8]~5 (
	.dataa(!\internal_counter[8]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\counter_snapshot[8]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \counter_snapshot[8]~5 .extended_lut = "off";
defparam \counter_snapshot[8]~5 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \counter_snapshot[8]~5 .shared_arith = "off";

dffeas \counter_snapshot[8] (
	.clk(clk),
	.d(\counter_snapshot[8]~5_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[8]~q ),
	.prn(vcc));
defparam \counter_snapshot[8] .is_wysiwyg = "true";
defparam \counter_snapshot[8] .power_up = "low";

dffeas \counter_snapshot[24] (
	.clk(clk),
	.d(\internal_counter[24]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[24]~q ),
	.prn(vcc));
defparam \counter_snapshot[24] .is_wysiwyg = "true";
defparam \counter_snapshot[24] .power_up = "low";

cyclonev_lcell_comb \read_mux_out[8]~28 (
	.dataa(!A_mem_baddr_2),
	.datab(!A_mem_baddr_3),
	.datac(!\counter_snapshot[8]~q ),
	.datad(!\counter_snapshot[24]~q ),
	.datae(!A_mem_baddr_4),
	.dataf(!\period_h_register[8]~q ),
	.datag(!\period_l_register[8]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[8]~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[8]~28 .extended_lut = "on";
defparam \read_mux_out[8]~28 .lut_mask = 64'hFF6FFFF6FF6FFFF6;
defparam \read_mux_out[8]~28 .shared_arith = "off";

cyclonev_lcell_comb \counter_snapshot[9]~6 (
	.dataa(!\internal_counter[9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\counter_snapshot[9]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \counter_snapshot[9]~6 .extended_lut = "off";
defparam \counter_snapshot[9]~6 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \counter_snapshot[9]~6 .shared_arith = "off";

dffeas \counter_snapshot[9] (
	.clk(clk),
	.d(\counter_snapshot[9]~6_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[9]~q ),
	.prn(vcc));
defparam \counter_snapshot[9] .is_wysiwyg = "true";
defparam \counter_snapshot[9] .power_up = "low";

dffeas \counter_snapshot[25] (
	.clk(clk),
	.d(\internal_counter[25]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[25]~q ),
	.prn(vcc));
defparam \counter_snapshot[25] .is_wysiwyg = "true";
defparam \counter_snapshot[25] .power_up = "low";

cyclonev_lcell_comb \read_mux_out[9]~24 (
	.dataa(!A_mem_baddr_2),
	.datab(!A_mem_baddr_3),
	.datac(!\counter_snapshot[9]~q ),
	.datad(!\counter_snapshot[25]~q ),
	.datae(!A_mem_baddr_4),
	.dataf(!\period_h_register[9]~q ),
	.datag(!\period_l_register[9]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[9]~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[9]~24 .extended_lut = "on";
defparam \read_mux_out[9]~24 .lut_mask = 64'hFF6FFFF6FF6FFFF6;
defparam \read_mux_out[9]~24 .shared_arith = "off";

cyclonev_lcell_comb \counter_snapshot[15]~7 (
	.dataa(!\internal_counter[15]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\counter_snapshot[15]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \counter_snapshot[15]~7 .extended_lut = "off";
defparam \counter_snapshot[15]~7 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \counter_snapshot[15]~7 .shared_arith = "off";

dffeas \counter_snapshot[15] (
	.clk(clk),
	.d(\counter_snapshot[15]~7_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[15]~q ),
	.prn(vcc));
defparam \counter_snapshot[15] .is_wysiwyg = "true";
defparam \counter_snapshot[15] .power_up = "low";

dffeas \counter_snapshot[31] (
	.clk(clk),
	.d(\internal_counter[31]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[31]~q ),
	.prn(vcc));
defparam \counter_snapshot[31] .is_wysiwyg = "true";
defparam \counter_snapshot[31] .power_up = "low";

cyclonev_lcell_comb \read_mux_out[15]~20 (
	.dataa(!A_mem_baddr_2),
	.datab(!A_mem_baddr_3),
	.datac(!\counter_snapshot[15]~q ),
	.datad(!\counter_snapshot[31]~q ),
	.datae(!A_mem_baddr_4),
	.dataf(!\period_h_register[15]~q ),
	.datag(!\period_l_register[15]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[15]~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[15]~20 .extended_lut = "on";
defparam \read_mux_out[15]~20 .lut_mask = 64'hFF6FFFF6FF6FFFF6;
defparam \read_mux_out[15]~20 .shared_arith = "off";

dffeas \counter_snapshot[12] (
	.clk(clk),
	.d(\internal_counter[12]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[12]~q ),
	.prn(vcc));
defparam \counter_snapshot[12] .is_wysiwyg = "true";
defparam \counter_snapshot[12] .power_up = "low";

dffeas \counter_snapshot[28] (
	.clk(clk),
	.d(\internal_counter[28]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[28]~q ),
	.prn(vcc));
defparam \counter_snapshot[28] .is_wysiwyg = "true";
defparam \counter_snapshot[28] .power_up = "low";

cyclonev_lcell_comb \read_mux_out[12]~16 (
	.dataa(!A_mem_baddr_2),
	.datab(!A_mem_baddr_3),
	.datac(!\counter_snapshot[12]~q ),
	.datad(!\counter_snapshot[28]~q ),
	.datae(!A_mem_baddr_4),
	.dataf(!\period_h_register[12]~q ),
	.datag(!\period_l_register[12]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[12]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[12]~16 .extended_lut = "on";
defparam \read_mux_out[12]~16 .lut_mask = 64'hFFF6FFF6FFF6FFF6;
defparam \read_mux_out[12]~16 .shared_arith = "off";

dffeas \counter_snapshot[13] (
	.clk(clk),
	.d(\internal_counter[13]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[13]~q ),
	.prn(vcc));
defparam \counter_snapshot[13] .is_wysiwyg = "true";
defparam \counter_snapshot[13] .power_up = "low";

dffeas \counter_snapshot[29] (
	.clk(clk),
	.d(\internal_counter[29]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[29]~q ),
	.prn(vcc));
defparam \counter_snapshot[29] .is_wysiwyg = "true";
defparam \counter_snapshot[29] .power_up = "low";

cyclonev_lcell_comb \read_mux_out[13]~12 (
	.dataa(!A_mem_baddr_2),
	.datab(!A_mem_baddr_3),
	.datac(!\counter_snapshot[13]~q ),
	.datad(!\counter_snapshot[29]~q ),
	.datae(!A_mem_baddr_4),
	.dataf(!\period_h_register[13]~q ),
	.datag(!\period_l_register[13]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[13]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[13]~12 .extended_lut = "on";
defparam \read_mux_out[13]~12 .lut_mask = 64'hFFF6FFF6FFF6FFF6;
defparam \read_mux_out[13]~12 .shared_arith = "off";

cyclonev_lcell_comb \counter_snapshot[14]~8 (
	.dataa(!\internal_counter[14]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\counter_snapshot[14]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \counter_snapshot[14]~8 .extended_lut = "off";
defparam \counter_snapshot[14]~8 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \counter_snapshot[14]~8 .shared_arith = "off";

dffeas \counter_snapshot[14] (
	.clk(clk),
	.d(\counter_snapshot[14]~8_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[14]~q ),
	.prn(vcc));
defparam \counter_snapshot[14] .is_wysiwyg = "true";
defparam \counter_snapshot[14] .power_up = "low";

dffeas \counter_snapshot[30] (
	.clk(clk),
	.d(\internal_counter[30]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[30]~q ),
	.prn(vcc));
defparam \counter_snapshot[30] .is_wysiwyg = "true";
defparam \counter_snapshot[30] .power_up = "low";

cyclonev_lcell_comb \read_mux_out[14]~8 (
	.dataa(!A_mem_baddr_2),
	.datab(!A_mem_baddr_3),
	.datac(!\counter_snapshot[14]~q ),
	.datad(!\counter_snapshot[30]~q ),
	.datae(!A_mem_baddr_4),
	.dataf(!\period_h_register[14]~q ),
	.datag(!\period_l_register[14]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[14]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[14]~8 .extended_lut = "on";
defparam \read_mux_out[14]~8 .lut_mask = 64'hFF6FFFF6FF6FFFF6;
defparam \read_mux_out[14]~8 .shared_arith = "off";

endmodule

module first_nios2_system_first_nios2_system_tenOut1 (
	readdata_0,
	readdata_1,
	readdata_2,
	readdata_3,
	Equal0,
	r_sync_rst,
	clk_clk,
	tenout1_external_connection_export_0,
	tenout1_external_connection_export_1,
	tenout1_external_connection_export_2,
	tenout1_external_connection_export_3)/* synthesis synthesis_greybox=1 */;
output 	readdata_0;
output 	readdata_1;
output 	readdata_2;
output 	readdata_3;
input 	Equal0;
input 	r_sync_rst;
input 	clk_clk;
input 	tenout1_external_connection_export_0;
input 	tenout1_external_connection_export_1;
input 	tenout1_external_connection_export_2;
input 	tenout1_external_connection_export_3;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \readdata[0] (
	.clk(clk_clk),
	.d(tenout1_external_connection_export_0),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(Equal0),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_0),
	.prn(vcc));
defparam \readdata[0] .is_wysiwyg = "true";
defparam \readdata[0] .power_up = "low";

dffeas \readdata[1] (
	.clk(clk_clk),
	.d(tenout1_external_connection_export_1),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(Equal0),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_1),
	.prn(vcc));
defparam \readdata[1] .is_wysiwyg = "true";
defparam \readdata[1] .power_up = "low";

dffeas \readdata[2] (
	.clk(clk_clk),
	.d(tenout1_external_connection_export_2),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(Equal0),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_2),
	.prn(vcc));
defparam \readdata[2] .is_wysiwyg = "true";
defparam \readdata[2] .power_up = "low";

dffeas \readdata[3] (
	.clk(clk_clk),
	.d(tenout1_external_connection_export_3),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(Equal0),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_3),
	.prn(vcc));
defparam \readdata[3] .is_wysiwyg = "true";
defparam \readdata[3] .power_up = "low";

endmodule

module first_nios2_system_first_nios2_system_tenOut1_1 (
	readdata_0,
	readdata_1,
	readdata_2,
	readdata_3,
	Equal0,
	r_sync_rst,
	clk_clk,
	tenout2_external_connection_export_0,
	tenout2_external_connection_export_1,
	tenout2_external_connection_export_2,
	tenout2_external_connection_export_3)/* synthesis synthesis_greybox=1 */;
output 	readdata_0;
output 	readdata_1;
output 	readdata_2;
output 	readdata_3;
input 	Equal0;
input 	r_sync_rst;
input 	clk_clk;
input 	tenout2_external_connection_export_0;
input 	tenout2_external_connection_export_1;
input 	tenout2_external_connection_export_2;
input 	tenout2_external_connection_export_3;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \readdata[0] (
	.clk(clk_clk),
	.d(tenout2_external_connection_export_0),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(Equal0),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_0),
	.prn(vcc));
defparam \readdata[0] .is_wysiwyg = "true";
defparam \readdata[0] .power_up = "low";

dffeas \readdata[1] (
	.clk(clk_clk),
	.d(tenout2_external_connection_export_1),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(Equal0),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_1),
	.prn(vcc));
defparam \readdata[1] .is_wysiwyg = "true";
defparam \readdata[1] .power_up = "low";

dffeas \readdata[2] (
	.clk(clk_clk),
	.d(tenout2_external_connection_export_2),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(Equal0),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_2),
	.prn(vcc));
defparam \readdata[2] .is_wysiwyg = "true";
defparam \readdata[2] .power_up = "low";

dffeas \readdata[3] (
	.clk(clk_clk),
	.d(tenout2_external_connection_export_3),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(Equal0),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_3),
	.prn(vcc));
defparam \readdata[3] .is_wysiwyg = "true";
defparam \readdata[3] .power_up = "low";

endmodule
